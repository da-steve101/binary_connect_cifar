`timescale 1 ns/1 ps

module aws_vgg_testbench;

wire [47:0] airplane4_image [1023:0] = { 48'h1100120014, 48'h1100130014, 48'h1200130015, 48'h1200130015, 48'h1300140015, 48'h1200130015, 48'h1200130015, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1400150016, 48'h1400150016, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1200130015, 48'h1200130015, 48'h1100120014, 48'h1100120014, 48'h1100120014, 48'h1100110014, 48'h1000110014, 48'h1000100013, 48'hf000f0012, 48'he000f0011, 48'he000e0011, 48'hd000e0011, 48'he000f0011, 48'h1100120014, 48'h1100130014, 48'h1200130015, 48'h1300130015, 48'h1300140015, 48'hf00100011, 48'hd000e000f, 48'h1200130015, 48'h1400150016, 48'h1300140015, 48'h1300140016, 48'h1300140015, 48'h1300140015, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1300140015, 48'h1200130015, 48'h1200130015, 48'h1100120014, 48'h1100120014, 48'h1100110014, 48'h1000110014, 48'h1000100013, 48'hf00100013, 48'hf00100013, 48'he000f0012, 48'he000f0011, 48'hd000e0011, 48'he000f0011, 48'h1100120014, 48'h1100130014, 48'h1100130014, 48'h1300140016, 48'h9000b000f, 48'h600090009, 48'h500050008, 48'h600060009, 48'h1000120013, 48'h1400150016, 48'h1300140015, 48'h1300140015, 48'h1200140015, 48'h1300150015, 48'h1300140015, 48'h1300140015, 48'h1300140015, 48'h1300140015, 48'h1200130015, 48'h1200130015, 48'h1100130015, 48'h1100120014, 48'h1100120014, 48'h1100110014, 48'h1000110014, 48'hf00100013, 48'hf00100013, 48'hf00100013, 48'he000e0012, 48'hd000e0011, 48'hd000e0010, 48'he000f0012, 48'h1100120014, 48'h1100130014, 48'h1100120014, 48'h1200140015, 48'hfffe00020008, 48'hfff7fff90001, 48'h400040008, 48'h100020004, 48'h200040004, 48'hf000f0010, 48'h1400140015, 48'h1200140015, 48'h1100140014, 48'h1200150015, 48'h1000120013, 48'hf00100011, 48'h1200130015, 48'h1200130015, 48'h1100130014, 48'h1100120015, 48'h1100120015, 48'h1100120015, 48'h1100110014, 48'h1000110014, 48'h1000100013, 48'h1000100013, 48'hf00100013, 48'hf00100013, 48'he000e0013, 48'he000e0011, 48'hd000f0010, 48'he000f0011, 48'h1100120014, 48'h1100130014, 48'h1100120014, 48'h1100130014, 48'hc000d0013, 48'hfff5fff60005, 48'hfff4fff80000, 48'h60004, 48'hffff00020001, 48'hffff00000000, 48'hc000d000d, 48'h1300150015, 48'h1100130015, 48'h1200140016, 48'h1100120014, 48'h9000a000b, 48'h1300140016, 48'h1300140015, 48'h1200130015, 48'h1100120015, 48'h1100120015, 48'h1100110014, 48'h1000110014, 48'h1000100013, 48'hf00100013, 48'hf00100013, 48'hf00100013, 48'hf00100013, 48'he000f0012, 48'he000f0010, 48'hd000f000f, 48'he000f0011, 48'h1100120014, 48'h1100120014, 48'h1100120014, 48'h1100120014, 48'h1300130016, 48'h8000c0012, 48'hffedfff30000, 48'hfff4fffa0000, 48'h100030007, 48'h3, 48'hfffcfffdfffd, 48'h8000a000a, 48'h1400150017, 48'h1100110015, 48'h200030005, 48'hfff5fff7fff9, 48'h300040006, 48'h1000110013, 48'h1100120014, 48'h1100110014, 48'h1100120015, 48'h1100110014, 48'h1000110014, 48'h1000110014, 48'hf00100013, 48'hf00100013, 48'hf00100013, 48'hf00100013, 48'he000f0011, 48'hd000e0010, 48'hd000e0010, 48'he000f0010, 48'h1000110013, 48'h1100120014, 48'h1100120014, 48'h1100120014, 48'h1200120013, 48'h1000140013, 48'h4000a000f, 48'hfff0fff20003, 48'hfff6fff70003, 48'h20006, 48'hfffe00000001, 48'hfffbfffdfffd, 48'h200030004, 48'hfffbfffbffff, 48'hfff3fff3fff7, 48'hffebffebffee, 48'hfff9fff9fffc, 48'h1000100014, 48'hd000e0010, 48'he000f0012, 48'h1200130015, 48'h1100110014, 48'h1000110014, 48'h1000110014, 48'hf00100013, 48'hf00100013, 48'hf00100013, 48'he000f0012, 48'hd000e0010, 48'hd000e0011, 48'he000e0012, 48'hd000e0011, 48'h1000110013, 48'h1000110013, 48'h1000110013, 48'h1100120014, 48'h1200130014, 48'h1200120014, 48'h1100130014, 48'h400060010, 48'hffeefff10000, 48'hfff7fff80002, 48'hfffe00000003, 48'hfffe0000ffff, 48'hfff5fff6fff6, 48'hffedffedffef, 48'hfffafffafffd, 48'hfffafffbfffe, 48'hffffffff0003, 48'h1400140017, 48'hd000d0010, 48'ha000a000d, 48'h1000110013, 48'h1000110014, 48'h1000110014, 48'h1000110014, 48'h1000100013, 48'hf00100013, 48'hf00100013, 48'hf00100013, 48'he000e0011, 48'hb000b0011, 48'h900090010, 48'hc000c0011, 48'hf00110013, 48'h1000110013, 48'h1000110013, 48'h1000110013, 48'h1100110014, 48'h1300110015, 48'h1300110014, 48'h1100150015, 48'h3000c, 48'hfff1fff1fffb, 48'hfffeffff0003, 48'hfffcfffefffd, 48'hfff7fff8fff7, 48'hfff9fff9fffa, 48'hfffbfffcffff, 48'h70008000a, 48'h100020005, 48'hc000c000f, 48'hfff6fff6fffa, 48'hfff2fff2fff7, 48'h60007000a, 48'h1100130014, 48'h1000110013, 48'h1000110013, 48'hf00100013, 48'h1000100013, 48'hf00100013, 48'ha000a000e, 48'hfffefffe0003, 48'hffefffeffff7, 48'hffe7ffe7fff1, 48'h100010009, 48'hf00100011, 48'hf00110011, 48'hf00110012, 48'h1000120013, 48'h1000120013, 48'h1100120013, 48'h1100120013, 48'h1100120013, 48'h1100120014, 48'h300040007, 48'hfffcfffdffff, 48'hfffbfffdfffd, 48'hfffafffcfffb, 48'hfffeffffffff, 48'hfffafffbfffd, 48'hfffcfffdffff, 48'h100020004, 48'hfffafffbfffd, 48'hffeeffeefff3, 48'hffedffedfff2, 48'ha000b000d, 48'h1100120012, 48'h1000110012, 48'h1000110012, 48'hf00100012, 48'hb000c000f, 48'h10005, 48'hfff0fff1fff5, 48'hffe5ffe6ffe9, 48'hffd9ffdbffe1, 48'hffdeffe0ffe9, 48'h30005000b, 48'he000f000f, 48'he000f0010, 48'hf00100010, 48'hf00110011, 48'h1000110011, 48'h1000110011, 48'h1100110012, 48'h1100120012, 48'h1100110012, 48'hf00100011, 48'h10002, 48'hfff8fff9fffa, 48'hfffdfffffffe, 48'hfffeffffffff, 48'hffff00000002, 48'hfffcfffdffff, 48'hfff4fff5fff7, 48'hfff5fff6fff8, 48'h100010004, 48'hfff9fff9fffd, 48'h9000a000b, 48'h1000110012, 48'hf00100013, 48'he000f0011, 48'h200040006, 48'hfff3fff5fff8, 48'hffe9ffebffed, 48'hffe3ffe4ffe7, 48'hffdaffdcffdb, 48'hffd1ffd3ffd4, 48'hffeffff2fff5, 48'hc000e000f, 48'he000e000e, 48'he000e000e, 48'hf000f000f, 48'hf000f000f, 48'hf000f000f, 48'h1000100010, 48'h1100110011, 48'h1100110011, 48'h1000100011, 48'h1000110011, 48'hf00100010, 48'hffff00010000, 48'hfff9fffafffa, 48'hfffeffffffff, 48'h400050006, 48'hffff00000002, 48'hfffcfffdfffe, 48'hfff7fff7fff9, 48'h100020003, 48'h600070008, 48'h80009000b, 48'hf00100013, 48'h90009000e, 48'hfff7fff9fffc, 48'hffe5ffe9ffea, 48'hffe7ffeaffeb, 48'hfff1fff4fff5, 48'hfffcfffeffff, 48'hffeeffefffee, 48'hffedffeeffee, 48'h700070009, 48'ha000b000b, 48'he000d000d, 48'he000d000d, 48'hf000e000e, 48'hf000e000e, 48'hf000e000e, 48'hf000f000e, 48'h10000f000f, 48'h10000f000f, 48'h100010000f, 48'hf0010000f, 48'h100010000f, 48'hb000c000c, 48'hfffdfffefffd, 48'hfffafffbfffc, 48'hffff00000002, 48'hfffcfffdfffe, 48'hfffeffff0001, 48'hfffeffff0000, 48'hfff8fff9fff9, 48'h700080009, 48'ha000a000d, 48'h4, 48'hfff1fff2fff5, 48'hffe9ffecffee, 48'hfff3fff6fff8, 48'h300050006, 48'h9000a000b, 48'h400040004, 48'hfffcfffbfffc, 48'h800050007, 48'hb0008000a, 48'ha0008000a, 48'hd000b000a, 48'hd000b000b, 48'he000c000b, 48'he000c000c, 48'he000d000c, 48'he000d000d, 48'hf000e000d, 48'hf000e000d, 48'he000e000d, 48'he000f000c, 48'he000e000c, 48'he000e000e, 48'h900090009, 48'hfffafffafffc, 48'hfff9fff9fffb, 48'hfffeffff0000, 48'h100020004, 48'h300040006, 48'hfff8fff9fffa, 48'hfff7fff8fff9, 48'hfff2fff2fff6, 48'hffebffebffef, 48'hfff3fff4fff7, 48'h300040006, 48'hb000d000f, 48'h80009000a, 48'hffffffff, 48'hfffefffe, 48'h700050006, 48'hb00070008, 48'hb00060006, 48'hb00070007, 48'hb00090008, 48'hb000a0008, 48'hc000a0009, 48'hc000a000a, 48'hd000b000a, 48'hd000c000a, 48'hd000d000b, 48'hd000d000b, 48'hd000d000b, 48'hd000d000a, 48'hd000d000a, 48'hc000c000a, 48'hd000c000b, 48'h600060006, 48'hfffcfffdffff, 48'h200030004, 48'h100020004, 48'hfff5fff5fff7, 48'hffe9ffebffec, 48'hffe8ffe9ffeb, 48'hffe9ffe9ffed, 48'hfffafffafffe, 48'he00100011, 48'hd000e000e, 48'hffffffff0001, 48'hfffafff9fffa, 48'h500030000, 48'hb00080006, 48'ha00070005, 48'h900060003, 48'ha00050002, 48'ha00060004, 48'ha00080004, 48'hb00090005, 48'hb00090006, 48'hb00090007, 48'hd00090006, 48'hc000a0006, 48'hb000b0008, 48'hc000b0008, 48'hd000b0008, 48'he000a0008, 48'hd000a0008, 48'hc000a0008, 48'hb00090008, 48'h900080008, 48'hfff9fff9fffc, 48'hfff2fff3fff5, 48'hffe9ffebffed, 48'hffe6ffe7ffe9, 48'hffe9ffebffec, 48'hfff9fffafffc, 48'h80007000b, 48'hc000c000f, 48'h200050006, 48'hfffcfffffffd, 48'hfffdfffcffff, 48'hfffbfffcfffe, 48'h40004ffff, 48'h900050002, 48'h800040001, 48'h800040000, 48'h700040000, 48'h800050001, 48'ha00060000, 48'hb00070001, 48'hb00070002, 48'hc00070003, 48'hc00070003, 48'hb00080004, 48'hb00090004, 48'hd00090004, 48'he00090004, 48'he00090004, 48'hc00080004, 48'ha00080005, 48'h900080008, 48'h600060007, 48'hffeffff0fff3, 48'hffdfffe0ffe3, 48'hffe3ffe5ffe8, 48'hfff2fff4fff8, 48'h300060009, 48'hc000e0010, 48'h80007000b, 48'hfffcfffbfffd, 48'hfff6fff8fff7, 48'h100040004, 48'hfff9fffbffff, 48'hffeaffebffed, 48'hfffcfffcfff8, 48'h800040000, 48'h70002fffe, 48'h70003fffd, 48'h60002fffc, 48'h70002fffd, 48'hb0004fffd, 48'ha0005ffff, 48'hb0005ffff, 48'hd0005fffe, 48'hb00050000, 48'hb00050000, 48'hb0006ffff, 48'he00070000, 48'he00060000, 48'hc00060000, 48'hb00070003, 48'h900060005, 48'h1, 48'hfff3fff4fff7, 48'hffe6ffe8ffeb, 48'hffe9ffebffee, 48'hfffe00010004, 48'he00100014, 48'ha000d000f, 48'hfffcfffd0000, 48'hfffafffafffd, 48'hfffefffeffff, 48'hfff8fff9fff7, 48'hfff9fffafffa, 48'hfff8fff8fff9, 48'hfff1ffefffed, 48'hfff9fff6fff1, 48'h70002fffa, 48'h60001fff9, 48'h60001fff9, 48'h60000fff8, 48'h60001fff9, 48'h80001fffb, 48'h70002fffe, 48'h80003fffd, 48'hb0004fffc, 48'hb0004fffd, 48'hb0004fffc, 48'hc0005fffb, 48'hb0005fffd, 48'hb0004ffff, 48'h900050001, 48'h40001fffe, 48'hfff8fff7fff7, 48'hffedffedffef, 48'hffeefff0fff2, 48'hfffbfffdfffe, 48'h9000a000b, 48'hd000d000d, 48'h500040002, 48'hfffafff9fff8, 48'hfffdfffcfffd, 48'h500060008, 48'h600070008, 48'hfffbfffcfffb, 48'hfff9fff8fff6, 48'hfffdfffbfff6, 48'h2fffdfff7, 48'hfff9fff3ffee, 48'h2fffcfff3, 48'h70000fff6, 48'h6fffffff4, 48'h6fffffff4, 48'h70000fff5, 48'h1fffcfff9, 48'h400000000, 48'h40001fffe, 48'h70001fffa, 48'ha0002fff9, 48'hb0003fff8, 48'hb0003fff7, 48'h90003fffb, 48'h40001fffd, 48'hfff8fff7fff7, 48'hffeeffedffee, 48'hffedffeeffef, 48'hfff5fff6fff9, 48'h500070009, 48'hb000d000e, 48'h500050003, 48'h2fffefff9, 48'h3fffefff5, 48'h1fffcfff5, 48'hfffefffbfff9, 48'h10001, 48'hfffe00000001, 48'hfffeffff0000, 48'hfffcfffafffb, 48'hfffcfffafff4, 48'h40000fffa, 48'hfffcfff8fff7, 48'hfff6fff3ffef, 48'h4fffdfff1, 48'h6fffefff1, 48'h5fffdfff0, 48'h6fffefff1, 48'h1fffafff5, 48'hfffffffafffc, 48'h200010004, 48'h40001fffe, 48'h6fffffff7, 48'h80001fff4, 48'ha0003fff7, 48'hfffefffafff4, 48'hffedffedffec, 48'hffe7ffe9ffeb, 48'hfff5fff7fff8, 48'h600080009, 48'hd000e000f, 48'h600060005, 48'hfffefffcfff7, 48'hfffffffbfff3, 48'h5fffefff3, 48'h9fffffff2, 48'h8fffefff2, 48'hfffffff9fff2, 48'hfffafff8fff6, 48'hfffcfffeffff, 48'hffff00010003, 48'hffffffff0002, 48'hfffafffafff9, 48'hfffffffefffb, 48'hfff6fff5fff8, 48'hffeaffebffe9, 48'hfffaffed, 48'h6fffdffee, 48'h4fffcffed, 48'h6fffdffed, 48'h9fffdfff0, 48'hfff8fff4, 48'hfffafffaffff, 48'h100020004, 48'h60002ffff, 48'h50000fff8, 48'hfffcfff8fff2, 48'hffeeffecffed, 48'hfff1fff3fff5, 48'h200030004, 48'ha000b000b, 48'h800080006, 48'h1fffffffa, 48'hfffffffafff2, 48'h5fffdfff0, 48'h8fffffff1, 48'h9ffffffef, 48'h8fffdffed, 48'h9fffeffed, 48'h8fffdfff0, 48'hfffafff2, 48'hfffdfffbfff9, 48'h2, 48'h200030004, 48'hfffdfffdfffe, 48'hfff8fff7fff5, 48'hfff9fff8fff5, 48'hfff6fff3ffeb, 48'hfffffff7ffe8, 48'h5fffbffeb, 48'h4fffaffe9, 48'h6fffaffe9, 48'h9fffcffeb, 48'h5fffcffee, 48'hfffafff7fff3, 48'hfffdfffcfffb, 48'h700040002, 48'hfffffffefffa, 48'hfff4fff4fff4, 48'hfffbfffafffd, 48'hfffffffffffe, 48'hfffffffd, 48'hfffdfff9, 48'hfffafff1, 48'h4fffbffee, 48'h8fffeffee, 48'h8fffeffee, 48'h8fffeffee, 48'h8fffdffed, 48'h8fffdffec, 48'h8fffdffec, 48'h8fffcffed, 48'h6fffbffed, 48'hfffffff8ffef, 48'hfffffffdfffa, 48'hfffe0000ffff, 48'hfff8fffcfff8, 48'hfffafff8fff8, 48'hfffcfff6ffed, 48'h2fff8ffe9, 48'h2fff6ffe6, 48'h5fff9ffe7, 48'h4fff8ffe6, 48'h5fff8ffe6, 48'h9fffaffe7, 48'h6fffcffe6, 48'h1fffaffeb, 48'hfffdfff7fff2, 48'hfffdfffafff9, 48'hfff5fff8fff8, 48'hfff3fff7fffa, 48'hffefffeffff2, 48'hfff4fff0ffeb, 48'hfffffff7ffec, 48'h4fffaffed, 48'h8fffcffec, 48'h9fffcffea, 48'h8fffcffea, 48'h7fffcffeb, 48'h7fffcffea, 48'h8fffbffe9, 48'h8fffbffe8, 48'h6fffaffe9, 48'h8fffaffe9, 48'hafffbffe6, 48'h6fff9ffe8, 48'hfffbfff5ffed, 48'hfff5fff7fff8, 48'hfff7fffcffff, 48'hfff8fff8fffb, 48'hfffcfff7ffec, 48'h4fff8ffe3, 48'h5fff8ffe5, 48'h4fff7ffe4, 48'h4fff6ffe2, 48'h5fff7ffe2, 48'h8fff9ffe5, 48'h6fffbffe1, 48'h6fffbffe4, 48'hfffcfff4ffeb, 48'hffebffe9ffe9, 48'hffe6ffe9ffe9, 48'hffe9ffebffee, 48'hfff2fff2fff4, 48'hfffbfff7fff0, 48'h7fffaffea, 48'hbfffcffe8, 48'hafffbffe6, 48'h6fffaffe7, 48'h5fff9ffe8, 48'h6fffaffe8, 48'h7fffaffe7, 48'h8fffaffe6, 48'h8fffaffe5, 48'h6fff9ffe6, 48'h8fff9ffe5, 48'hafff9ffe2, 48'h8fff9ffe3, 48'h1fff7ffe7, 48'hfff3ffefffed, 48'hfff1fff1fffc, 48'hfff3fff7fffa, 48'hfff8fff7fff2, 48'hfffefff6ffe4, 48'h3fff7ffe1, 48'h3fff5ffe1, 48'h3fff5ffe0, 48'h5fff6ffe0, 48'h5fff7ffe3, 48'h5fff8ffe1, 48'h8fff9ffe1, 48'hfffbfff2ffe5, 48'hffe1ffe1ffe2, 48'hffe0ffe2ffe2, 48'hffeeffedffeb, 48'hfffbfff9fffa, 48'hfffefffcfff8, 48'h1fff8ffeb, 48'h6fff8ffe6, 48'h9fff9ffe3, 48'h8fff9ffe3, 48'h5fff8ffe4, 48'h5fff8ffe4, 48'h6fff8ffe3, 48'h6fff8ffe3, 48'h7fff8ffe2, 48'h6fff8ffe2, 48'h6fff8ffe2, 48'h6fff7ffe1, 48'h6fff7ffe1, 48'h5fff7ffe1, 48'hfffffff3ffe6, 48'hfff3ffeeffee, 48'hffeeffeffff6, 48'hfff3fff4fff8, 48'hfffbfff5ffee, 48'hfffffff4ffdf, 48'h1fff4ffde, 48'h1fff4ffdd, 48'h3fff5ffdd, 48'h3fff5ffe1, 48'h4fff6ffe0, 48'h8fff7ffde, 48'hfff8fff0ffe3, 48'hffe0ffe1ffe3, 48'hffe7ffe7ffe4, 48'hfff7fff1ffe8, 48'hfffafff3ffec, 48'hfffdfff9fff4, 48'hfffbfff4, 48'h1fff6ffe7, 48'h7fff7ffe1, 48'h9fff8ffdf, 48'h7fff7ffe0, 48'h5fff7ffe1, 48'h5fff6ffe0, 48'h6fff6ffe0, 48'h6fff6ffe0, 48'h6fff6ffdf, 48'h5fff6ffdf, 48'h4fff5ffe0, 48'h4fff5ffdf, 48'h6fff5ffdd, 48'h6fff5ffdd, 48'hfffdfff4ffe0, 48'hfff0ffecffed, 48'hfff1ffeffff8, 48'hfffafff7fffa, 48'hfffefff4ffe4, 48'hfffffff2ffdd, 48'h1fff3ffdc, 48'h3fff4ffdb, 48'h3fff4ffdf, 48'h4fff5ffdd, 48'h7fff6ffdb, 48'hfff4ffedffe3, 48'hffdfffe1ffe3, 48'hffedffe9ffe2, 48'h2fff4ffe2, 48'h3fff4ffe0, 48'hfffffff4ffe5, 48'hfff7ffec, 48'h2fff5ffe4, 48'h6fff5ffde, 48'h6fff6ffdd, 48'h5fff5ffde, 48'h6fff5ffde, 48'h6fff5ffde, 48'h5fff5ffdd, 48'h5fff5ffdd, 48'h5fff4ffdd, 48'h5fff4ffdd, 48'h5fff4ffdd, 48'h5fff4ffdd, 48'h5fff4ffdd, 48'h5fff4ffdc, 48'h2fff5ffda, 48'hfffafff1ffe1, 48'hfff3ffecffed, 48'hfff8fff4fff3, 48'hfffefff4ffe7, 48'hfffefff1ffdd, 48'h2fff2ffda, 48'h4fff2ffda, 48'h3fff3ffdd, 48'h3fff3ffdb, 48'h5fff4ffda, 48'hfff4ffecffe0, 48'hffe6ffe4ffe0, 48'hfff4ffedffe1, 48'h4fff4ffdd, 48'h6fff5ffdc, 48'h1fff3ffdf, 48'hfff3ffe1, 48'h4fff4ffde, 48'h6fff4ffdc, 48'h4fff4ffdc, 48'h3fff4ffdd, 48'h5fff4ffdc, 48'h5fff4ffdc, 48'h4fff3ffdb, 48'h4fff3ffdb, 48'h4fff3ffdb, 48'h4fff3ffdc, 48'h4fff3ffdb, 48'h4fff3ffdb, 48'h4fff3ffdb, 48'h6fff2ffdc, 48'h5fff3ffd8, 48'h2fff2ffdb, 48'hfffdffefffe1, 48'hfffcfff1ffdf, 48'hfffefff1ffdd, 48'hfffffff1ffda, 48'h1fff1ffd8, 48'h2fff1ffd8, 48'h3fff2ffdb, 48'h4fff2ffda, 48'h5fff3ffda, 48'hfff9ffedffdd, 48'hfff2ffebffde, 48'hfffdfff2ffdf, 48'h5fff4ffda, 48'h6fff4ffd8, 48'h4fff3ffdb, 48'h4fff3ffdb, 48'h6fff3ffda, 48'h6fff4ffda, 48'h4fff3ffdb, 48'h3fff3ffdc, 48'h4fff3ffdb, 48'h4fff3ffdb, 48'h4fff2ffda, 48'h4fff2ffda, 48'h4fff2ffda, 48'h4fff3ffda, 48'h4fff2ffda, 48'h4fff2ffda, 48'h4fff2ffda, 48'h4fff1ffda, 48'h5fff2ffd7, 48'h4fff2ffd7, 48'h4fff1ffda, 48'h4fff1ffd7, 48'h2fff1ffd8, 48'hfff0ffd7, 48'hfff0ffd6, 48'hfff0ffd7, 48'h3fff1ffda, 48'h4fff1ffda, 48'h4fff1ffda, 48'hfff1ffdc, 48'hfffdfff1ffdd, 48'h1fff2ffdb, 48'h5fff3ffd8, 48'h6fff3ffd8, 48'h5fff3ffd8, 48'h5fff3ffd8, 48'h6fff3ffd8, 48'h5fff3ffd8, 48'h4fff2ffd9, 48'h3fff2ffda, 48'h4fff2ffd9, 48'h4fff2ffd9, 48'h4fff2ffd9, 48'h4fff2ffd9, 48'h4fff2ffd9, 48'h3fff2ffd8, 48'h3fff1ffd8, 48'h3fff1ffd8, 48'h3fff1ffd8, 48'h2fff1ffd7, 48'h1fff1ffd6, 48'h2fff1ffd8, 48'h3ffefffd9, 48'h3ffeeffd9, 48'h2ffefffd6, 48'hffefffd5, 48'hffffffeeffd5, 48'hffffffeeffd6, 48'h3fff0ffd7, 48'h4ffefffd8, 48'h2ffefffda, 48'h2fff1ffd9, 48'h2fff1ffd9, 48'h2fff1ffd9, 48'h4fff1ffd8, 48'h4fff2ffd8, 48'h4fff2ffd8, 48'h4fff2ffd7, 48'h4fff2ffd7, 48'h4fff1ffd8, 48'h4fff1ffd8, 48'h4fff1ffd8, 48'h3fff1ffd8, 48'h3fff1ffd8, 48'h3fff1ffd7, 48'h3fff1ffd7, 48'h3fff1ffd7, 48'h2fff0ffd7, 48'h2fff0ffd7, 48'h2fff0ffd7, 48'h2fff0ffd7, 48'h1fff0ffd6, 48'hffefffd7, 48'hffefffd7, 48'hffeeffd7, 48'hffedffd7, 48'hffedffd6, 48'hffffffedffd5, 48'hfffdffecffd5, 48'hffedffd5};

   wire [127:0] airplane4_mp_2_image [1023:0] = { 128'h6001e002700060005003400230006, 128'he000d00010000001800040008, 128'h17000000050018000600000007, 128'he0017001a00080000000a0010001e, 128'h180005001100130005000d00020000, 128'he0000001000010002001e001a0013, 128'hc00020028000b0016000300060017, 128'h12001d00000014000e00000008001a, 128'h8000b0000001e00060014001f0015, 128'h180000000500180009000c0014, 128'h11000000070000000000240007000d, 128'h400000029001700000013000a0013, 128'h120002000000060022000d00060010, 128'h18000000060003000c000700000000, 128'ha0012001200070000000a0011000a, 128'h60009000700100000000000030013, 128'h2500000013003700200008, 128'h13000000000002001000000000, 128'h16000000130014, 128'hd00080028001600040015001a0025, 128'h3e001b002b0003001e000c00000008, 128'h330005000c00070000000000160000, 128'ha001200120000001e0000000d000d, 128'h1a0018000000010002000000000026, 128'h1b0020000a000b00070011004d0000, 128'hd000f000800000018000e00040023, 128'h90006000c0000000b001300040019, 128'hb0000001c004d000b0000000d0000, 128'h220000002b0000002c000000130010, 128'h31000000000001001c000000000000, 128'h8000300000007000000180001000b, 128'hf000300040007000c00000004000e, 128'h3000000022000800000007, 128'h13000000000000, 128'h110000001c002300030000002a, 128'h800000022000a0003000000000014, 128'h30001a002700000026000000000007, 128'h2e0019001d00010000000e00000000, 128'h110000001c0002000d00000000, 128'h12000000000000001300000001002a, 128'h2300060000000000050010004a0000, 128'h13000e0000001d000000050014, 128'h1d0000001d002a00190005, 128'hb00310000000000140005, 128'h18000000380000002a0000001b001d, 128'h1c0000000d00110004000000000000, 128'h500100000001b0000000800080000, 128'h600000000001b, 128'h4000050000000400000000, 128'h3000e000b001c000600000000, 128'hb00000003000f002d00100011002b, 128'he0003002b0000000000000010001f, 128'he0000001100070009000000000000, 128'h420015002300000000001900060003, 128'he00120003000c000e00000009, 128'h18000d000000010011000000000011, 128'h20000d00000012000c001500150000, 128'h11000c0008001e000000040000, 128'h20000001200000007001900180000, 128'hb001900160000000f00140012, 128'h130000000e00000022000000140026, 128'h2100010000001f000d000a0005000d, 128'hb0000000a0000002300150000, 128'h2000000020006000000000016, 128'h1c00000000000000040001, 128'h1200120000000900000000, 128'hf0000000a002000120001001c, 128'hd0000002700000002000500090021, 128'h80000000a00000012000000000000, 128'h3800000019000100000017000f0000, 128'h3000e00000006000d000a00000003, 128'h16001300000003000b00000001000a, 128'h2a00120000000a000a001400030000, 128'h9001c0003000e00210000000a0009, 128'he0002002100000009001b00260002, 128'h12000f000e000000130014000e, 128'h180001002200000023000000150017, 128'h210004000d00000009000500030000, 128'he0021000000070000002200210000, 128'hb000d000000000022, 128'h1000500000000000000070004, 128'h800110004000e000e0000, 128'he000100080022001700000000, 128'ha000100100000000000020000000c, 128'hf0000000b000000000000, 128'h170000001a0000000000170011000e, 128'h500100007000b000e000d00000001, 128'h1200000006000e000000000008, 128'h200000000000170007001700050001, 128'h1e00000000001f000400090014, 128'h60000001900000008000600240000, 128'h7000000060008000000120018000b, 128'hd0000000c0000001700020012000b, 128'h18000000000000000e0005000a0000, 128'h30000000a00070000000800250000, 128'h4001100000000000b, 128'h4000b00000000000300070001, 128'h500110007000d000e0000, 128'hf000100070021001700000000, 128'ha0005000d0000000000020000000a, 128'he00000000000300030000, 128'h4000000220000000000180012000f, 128'h120003000a000d000c00000005, 128'h1200000004000900000000000a, 128'h220000000000160000001800050000, 128'h1e00030000001a000500090013, 128'ha00000006000000080007001f0000, 128'h7000000050008000000130018000b, 128'h4000100000001001300010012000d, 128'h16000000000000000f0000000a0000, 128'h20000000e00060000000300260000, 128'h10005001200000000000d, 128'h1d001500020000000f00160003, 128'h80000000f0014000d001600150006, 128'h3000a001c000a0023001700010004, 128'he00080011000c000000040004000d, 128'h80003001100090000000c00130000, 128'h15000c001e00000000001c0010000d, 128'h2000c002100080011000c00000013, 128'h2000f00000006000700080003000d, 128'h1a000d0001001e000300190002000c, 128'h28000500000020000b000b0014, 128'h8000d0006000200080003001a0006, 128'h90000000c0006000b000c00160015, 128'h500090005000b0018000b00100022, 128'h1500000000000d000a000700130018, 128'h600000007000b0000001800260004, 128'h500050000000c000200170004, 128'h40033000400000000002200080023, 128'h3000b00080000001a00040000, 128'h2a0000000a0011001300000000, 128'hd0001000000000006000000000000, 128'ha0004000700000013000e00000000, 128'h700000002000000110006000f001c, 128'h250006000d000000170000, 128'h2000e00000015000f000400190030, 128'h200010000000e00120000, 128'h1f000000000007000000080000, 128'h130000000f00000014001600300000, 128'hf0000000d00100000001700000003, 128'h20001000f00150009000f0000, 128'h18000000130000000d000000220004, 128'h30009001e0014000000160000000c, 128'he001e001f00050012001a, 128'h3f00000000000d004e00000019, 128'hd002300000000, 128'hf000000000000001b00000009, 128'h270000000000000000000000040000, 128'h3700020012000c001a000000000013, 128'h500000004000000080000000b0028, 128'he0000002200200000001100250000, 128'h5000000000000000000000017004c, 128'h100000000000000014000a00540000, 128'h260000001c, 128'he0000000800000049000200080005, 128'h500000018003a000d000000000000, 128'h1b0000000000000009000000000000, 128'h140000000000000010000000100005, 128'h1c00370000000600000012, 128'h1a0000001d0024001a000000000019, 128'h14000000320000002d003d00000000, 128'h10000000000021000600000000, 128'h1e0000000f001800000000000d000a, 128'h3800000000000c00000000000d0000, 128'h340012000400070017000000110022, 128'h250011001500000000000000000014, 128'h80000000300370000000b00220000, 128'hf000000000000001f0007000a0025, 128'h900000000001100160005005e0000, 128'h25000600000000002100000029, 128'h2400030036000000000003, 128'h1b001f000e000000010000, 128'h120000001a002a001d000000090000, 128'h8000a001b0000000000080014, 128'h17000000320000000000000000, 128'h110000000b00000000000000000000, 128'h430003000f0012000b0000, 128'hc000f00000000001d00040000000e, 128'hf0000000200140000000000350020, 128'h7001a001c00000006002a0011, 128'h26001c000000090006000b0011000b, 128'h2f001d000000080000000000160000, 128'h2001d0007000000140000000b0000, 128'h1a000000100003001e000e000c000d, 128'he000f000000260006001300190017, 128'h2d002100050000001200010000000f, 128'h2001e00000000000400000006, 128'h27001d0006002600000000000b, 128'h10004001c000a000300000014, 128'h380000002a001a0000000c0015, 128'he000c000200100000000900000014, 128'h30020002000010000000000000014, 128'ha003e0000000a001300140000, 128'hf002600120016000a000000060021, 128'h1400000000003e0029, 128'h80002001a001e0013000000150004, 128'h23000a0000000f0024000700000017, 128'h310016001a000c000b00150004000a, 128'ha0000000f0007000000030000, 128'h270000000d0003000000000000000d, 128'h240013000a0000001800020011001d, 128'hf00000000000f00100001000a0000, 128'h6000900330004000b002c00000004, 128'h2c001c0009001a000000000013, 128'hd00090025000e0020000000000010, 128'hd002c0013000d0000000300000008, 128'hf0028000000000001000700000022, 128'h1b000e001300170000000000050038, 128'h3300050004000000000004, 128'h2000e001a0024000000000000, 128'h170009000000230028, 128'h1c0005001100000013000000060000, 128'hb0000000000000022000000000000, 128'h2d0004001000000007001c00040009, 128'hb0000000c0000000f00000000, 128'h9000000160007001900000000000f, 128'h2200000004000100030000000f0000, 128'h30001000000000017000000000000, 128'h7000c003f0000000b0022001b0000, 128'h1b00000000000500000000000e, 128'h15000700290000001c00030011000b, 128'h60014001800060000000000040000, 128'h50022000a00000000002500000000, 128'h8000000160002000000040034, 128'h3900170000000300000000, 128'ha00170021000000000001, 128'h11000000000007001d000800000016, 128'h180011001800000005000200270015, 128'h1a0000000000000000, 128'h1e00030016000000000010000d0025, 128'h80028000d0004001b0000001b, 128'h5000f000e0000001800000000000a, 128'h1c00230002001400020000000c0000, 128'h100020000000b000000030000, 128'h1400000007000000110000, 128'hb00000000000000020000, 128'h3000000010000000e0000000e0010, 128'h3000400000029000d000000360002, 128'ha001200000000003c00000000, 128'h1e0000000800140017000e0001, 128'h1000a002e00100000000c00000001, 128'h240003001d0008000000020000000b, 128'ha00000016001600180000001e0029, 128'h130021003300130002002000300028, 128'h110000000000150002000600100009, 128'h30000f001a000000030007000f0008, 128'h7002900110017000d00000018, 128'ha0007000f00000000000000000009, 128'h21003e000b00140000000000000004, 128'h3c001a000c000b001e0000001a0000, 128'h130009001c0001000c000c00070007, 128'h2d002e00100000000000000009, 128'hd000600110000001f0001000d002b, 128'h2b000c0000001e00090000002a0024, 128'h3e001900020001000c004300000000, 128'h1e0000000300000014002a0026, 128'h600160005000000010005000e001b, 128'h3000a000d0000000000020000, 128'h2500000008000b000000060000, 128'hf0000000000070012000000000000, 128'h90000001b000b00000000, 128'he0005000d00100008001f, 128'h80000000700050000, 128'hf00130000000e0009000000050018, 128'ha000000060000000b000000060000, 128'h1100000000000b0000000c0000, 128'h7000000150000000c001b002f0000, 128'hd0000001000000004001300000008, 128'h2000e000f0015000d00160000, 128'h110000001a000a000a000000210000, 128'h1b002000090006001c00060000, 128'h160000000000190019000e000b0014, 128'h3e000000000000001f00000024, 128'h1d00000000, 128'h13000000000008001600070000, 128'h110000000000000000000000000000, 128'h60000000500000000, 128'h6000000120000000b0024, 128'h1e000000000006001b0000, 128'h5000000000001000000190029, 128'h90000000000070000000700000000, 128'h3000000000000000000000000, 128'hb000000120000002f0000002d0000, 128'h500020000, 128'h20000000900190000001b0000, 128'h100000000000300140000002d0014, 128'h1c003d0000002400000000, 128'h300220019000b00030020, 128'hd003b00000000001a004a0000000f, 128'h14002000000000, 128'h130000001600000000001800000004, 128'h220000000000000000000000000000, 128'h30000001000060000000000070030, 128'h1b0000001400000006001a, 128'h13000b0026003f00000005001f0000, 128'h9000000000022001d001a001d, 128'h500000000000c0004000300230000, 128'h400000000000000240000000f, 128'hc000000130010002a000100170000, 128'h90000001700090000000000010000, 128'h16000000000003001b0000000d0000, 128'h30000000b001b, 128'h1400430000000e00000000, 128'h70009001300180005000000000016, 128'h160000000000110015001f00080008, 128'ha0000000000090010001e0006, 128'h1e000a00160000000b001300000004, 128'h2d0000000000000000000000080002, 128'h280031001800130000000000030020, 128'h50014000e0004000000000000001d, 128'he000e000400110009000500220012, 128'h20000000d00230022000c0014, 128'h230026000b, 128'h1e000800000000000800000003, 128'h6001600120003001c0000, 128'h14000000000012000e000000090000, 128'hd00000008002c001b0000001c0000, 128'h12000e0006000000080005, 128'h30000000c002c0000000c0000001b, 128'h40016001700000003000000000000, 128'h9000100090025001f0005, 128'h8002f000000000022000e00230027, 128'h1e000000020028000e000d0025001d, 128'hc000000290003000000150000, 128'h1c0024000b001d0004000000000025, 128'h1200170012000d0000000e0000003a, 128'h6000d000d0027000a00000019000e, 128'h1100000003000400050012000b000d, 128'h400000005001900250013, 128'h190017000b00000000000a00040002, 128'h60000000a000a001500080014, 128'hc001e000a0001002c000000000000, 128'h1000000210000001000060008, 128'h50014000500000000000600000019, 128'h60000000d000500000000001b, 128'h22000f001200000000000000000000, 128'h200000038001c00000000000b0000, 128'h190000002c00310000002b000d, 128'h3500000010002b0002000000220023, 128'ha0008000e001c000d00140000, 128'h1b0005000000140009000000010013, 128'h1b0006000e0000000d0032000a003e, 128'h300030000000200000026000c0008, 128'h1a0003004800010024000000030000, 128'h20000000d001d000000000023000c, 128'hb0000000000000019000000000000, 128'hc00000009001400070001, 128'h1f000e00050027000000140000, 128'h23002d0000001700000000, 128'hf00290018001e000000220000, 128'h2001b000f000000030000000b0009, 128'h1000360000000000000029000f0010, 128'h50034001d0000000000000000, 128'h22001c000000000001, 128'h30000001e0000000000000000000a, 128'h1b002c00060012002a00480006, 128'h1d0005001a002500000000000c0000, 128'h15000b0003000000000000001b000c, 128'h10000500200005002a00210000001a, 128'h44000000000000000d0000, 128'h80021000000390000000000000000, 128'h440009000f00000010000000000003, 128'h10000000000010000000000000014, 128'h100170018000e000000160000, 128'hd00000000000000090000, 128'h600000027003a001b00320010, 128'h1e0014001600000000002700000000, 128'h4f000000000000003100010002, 128'h25000000000005000900000000, 128'h210007000000090029000c002b000e, 128'h1a00180007000700000000001f000c, 128'h260012001b002a003100320002, 128'h190000002800080009000800160007, 128'h2400100000000d000d000000080000, 128'h12000d0005000f0023000000000000, 128'h9000d001000160001000a00200000, 128'hf001d000700180000000000000014, 128'h5e001a000700060012000b00110009, 128'h20000500090017000f0000000a0012, 128'h5002100220012002b000000000000, 128'h50011000000000000000000000000, 128'he000f000000060008001900110033, 128'h3d00000000000000180000001f0017, 128'h200025000300030021001a00030020, 128'h900010010000100040005000e0005, 128'h20007000e0000000000050000, 128'h1d00000009000b000000030006, 128'hb0000001100120016000000000006, 128'hf00020016000e00000000, 128'hf0008000700120005001d, 128'h4000200080000000e00000000, 128'h11000b0006000c0008000000000015, 128'h190004000b0004000b000000120000, 128'h800000000000a000600090000, 128'h70000001200000000001a00120010, 128'hc0007001400010008000a00050009, 128'h40017000700150013000c0000, 128'h130000001b001300090002000e0000, 128'h2100160001000d001a000d0000, 128'h190000000000100014000b00060010, 128'ha001900000000000000000015, 128'h110008000000000000, 128'h4001000010000000c00000000000c, 128'h110001001100000000000000000000, 128'h3000900000000, 128'h8000300110000000400000000001b, 128'h6000100020000000c00050000, 128'h9000000000015000000000013, 128'h210000000000050004000000000000, 128'h1000000000002000000000000, 128'h200000012000000150000002e0000, 128'h1000000070005, 128'h700040003000f0000001d0004, 128'h140009000200220000, 128'hd001900090000002700000000, 128'h17000d000f00050011, 128'h45000c00000002001c0000000e, 128'h70023000e00000004, 128'h2d000400120006002c000a0000000d, 128'h90021000600000000000000040000, 128'h120000000200000000, 128'h11000000190000001200000003003a, 128'h9000b001600180000000900090020, 128'h9000000000017000000130017, 128'h10000000000000003000000000000, 128'h6000000000000, 128'h8000000030000003a0000002a0000, 128'h4000000090000, 128'h400180013001a0013, 128'h1a000800000046001a, 128'h17002d0000002a00000000, 128'h8001b0017001400090022, 128'h16002c000700000000002800000000, 128'h90032001700000010, 128'h2a000000290010001c000000000019, 128'h210023000e00060000000000190000, 128'h300060000003e0000000000000021, 128'ha00000019000000160000000d0030, 128'h50000001b003c0000000b00050030, 128'h160032000000200000000b0011, 128'h7000e00000003000d00260000, 128'h14000000000000000f001400000006, 128'h10000002f000000000000, 128'hc0006000b00000007000000150000, 128'h140019000d00100002, 128'h60010001c00000000003c0023, 128'h1d00280002001b00000000, 128'h500230008000000000029001c0000, 128'ha0007000000210000000200020002, 128'h3b00030017000e, 128'h1f00000021000e000b000000000017, 128'h19000000130033001a000b0000, 128'h50000003c000000000003001d, 128'h800000000000000000030, 128'h20000000200140018003200000016, 128'h19003e00000006000000170000, 128'h23000400150000001200050000, 128'h110000002400070008000f00000000, 128'h240011000000130000, 128'hc000300150003000a000000320000, 128'h12000c0008000e0000, 128'ha000c0009001800000028000d, 128'h90002000000030007000500000000, 128'h2e002500000000002e00080000, 128'h150000002c0000000000140000, 128'h150030000000000000, 128'h1b0000001100000000000000000013, 128'h2e0017000000310028000e001e, 128'h21001600420005000000000000000d, 128'h1000100000000000000000006, 128'h300000000000c004800320000003f, 128'h12004600000015000100150000, 128'h22000000430000000900000000, 128'hb00240000000000000000, 128'h700100000000500000000, 128'hb000f00000000003f0000, 128'h20024001e0000000000010000, 128'h1e0001001a000000080000, 128'h9000a0000, 128'h4700000000000e000f00000000, 128'h240000000000020000, 128'h80018001e000000000000, 128'h2d002300000000000400000000, 128'hd002200240009000d002f00000004, 128'h30001c00530010000e00000000000c, 128'h160000000e0000000000000000000e, 128'h4001200050000003e002200000045, 128'h20000000a00050000000000110000, 128'h50003000000230000001a00000000, 128'h900020000001c0002000000070003, 128'hc000000000000000e001e, 128'h500230006000e001f0000, 128'h1a001c003c000d00000008000e0000, 128'h600000009000000280015000b0000, 128'h310000000000000000000f00120019, 128'h4200000000000d000000000003, 128'h160003000f0000001200060003, 128'h90000000b001c00250000002c0007, 128'hb0037000700000022000f0000000b, 128'hd000000140008001c00380000000a, 128'hd000500330006000f000000010001, 128'hc00030004001000000005001b, 128'h20001f00100005000b0009000b0029, 128'h28000300080016000000140019, 128'h80000001f0000001c0000000a, 128'h1000230025000000200008000a0009, 128'h1000000180000000500000025001a, 128'h60014000a001300060000, 128'h1d0015002800080000002500130018, 128'he0000001c000a0000001200030000, 128'h1d000000190000000b0029001e001b, 128'hf000000000000003e0000000a0003, 128'h2700000017000a0007002c0015000a, 128'h7000e00080000000900000008, 128'h30010000000080008000000040017, 128'h3200060019001c000b000000150011, 128'h17000b0010000e002d001900000003, 128'h120000001300080000000d00050012, 128'h9000b001b00210002001200050000, 128'h16000200080003000000000000001f, 128'h25000b000a000000180003001c0002, 128'h800000005000c000900060003000e, 128'h70014000f0009000c001c0003001f, 128'h200005001b00130003000c0009000a, 128'h200003001b000e00110000, 128'h14000700190015000f000200060002, 128'h1800130014001b001a00000002, 128'h1a00000000001c001c000700070010, 128'h3100000021000c0000000000000000, 128'h400000019001f000000000000, 128'h3c000000170007000b000000010015, 128'h220025001900070000000900100002, 128'h120019000400120000000500000009, 128'h22000e000200000000001d000d0027, 128'h3001300130000001000040026, 128'h7000b001800000018000000000007, 128'h1800060000000a0000000000220000, 128'h400020007001f000000000009, 128'h4000a0000000b0007000a001c, 128'h9000000080006, 128'h1e000d000e001c00070009, 128'h11002a0000000000280004, 128'hd001e00000000001b00000000, 128'h2b000000000000000f00000007, 128'he0000002700250000000000000000, 128'h21002a000000000000, 128'h370000001e0000000800000000001e, 128'h12002d00210002000f003700220000, 128'hc0000001f0000000000080002, 128'h20001100080000000000000014002d, 128'h30004000b002a00000031, 128'h13004300000011000000000000, 128'h7000a000000140000000000000000, 128'hf0000000a0001001d000000000001, 128'h110011000000150000, 128'h10002400000000001c0000, 128'hd000600000018000d0007, 128'h2b001e00000047000e, 128'h200008002d00000000003000000000, 128'h400000000000000030000f0007, 128'h1a000600320000000000060000, 128'h5003b000500000000, 128'hf0000002300000000000000000024, 128'h2e001a00040043002b000d0009, 128'he0006003800230000000000070000, 128'ha00000000000000000000, 128'h90010001100420028000a0028, 128'h20053000000000000001c0000, 128'h10015000d001f0000000400000000, 128'hf0000000900090002000000000002, 128'h1f00000000000b000a, 128'h13002a00000000002b0000, 128'ha0014000600000000000a0000, 128'h700130004002e0028, 128'h2b0000000500000010000000000000, 128'h37000b0000001e002b00110000, 128'h15000000350000000e000f0000, 128'h2a000000000000, 128'h4000d002600000000000000000000, 128'h3000130000004400260000000e, 128'h200020004c00120000000300000000, 128'hf0000000000000000000a, 128'h400000000004300310007002c, 128'h2003400000000000000200000, 128'hf0020000000350000001200000000, 128'h2100000009002c000000000000000d, 128'h5000000000000001f, 128'h1c001f000d000600290000, 128'h140020001200080000000000000000, 128'h1f000e00110000, 128'h80001000000000008001100130000, 128'h41001700000026000100000008, 128'hb000000020000001300120009, 128'h16000e002a000d00050000, 128'h2900000000001b000a00000005, 128'h180039000f00000000002500000000, 128'h2b00260050000d000000050000000f, 128'h4001000000000000000000020, 128'h16001300070000002000000010002f, 128'h3000c000a, 128'hb0000000000230000001d00000000, 128'h29001d000a00200000000000000000, 128'hb0013000d000000170004, 128'h200000000001d0021000100170000, 128'h29002b001600160000000000120000, 128'h110009000000000004000000000000, 128'h1b0000001100070000001100120010, 128'h160000000a0012000000000000, 128'h400070004000d0028001700000013, 128'h2000000001002a001800260012, 128'h11001d000000050018000600190016, 128'h80001000000240018000000000000, 128'h3000180025000d0029000b0000001e, 128'hc0016000600000000000000000025, 128'h22001a0017002300000001001a000b, 128'hf0000000000100005000000050018, 128'h90000000d00000015001300110000, 128'h210010000b00170000001000000007, 128'h800000016000200280008000b0027, 128'hc000400280028000000000000, 128'hf0013002e001f0003000e00000000, 128'h18000a001f00000000000a00000011, 128'h1a000a0010000d001400000000001b, 128'h210000000000040000000000000010, 128'h160000000c0009001100020000000b, 128'h90024000e00100007000000000000, 128'h70018000b0000001a0000001f0010, 128'h17000000090014001f000000020008, 128'h1b000000130008002a000c00070010, 128'h170005000000080003001300000014, 128'h3000b00130003000b000a0004, 128'h80009000d000a0015000000020019, 128'hf0001000b00100017000700110008, 128'hb0024000a000f002200030000000b, 128'h2900000001001200170023, 128'h2a00050006000000000000000c, 128'h1e0003003b0013001f001f00100016, 128'hd000d003000170002000400050000, 128'he0028002400010011002f00050009, 128'hc00030002000000050009000d0014, 128'h1e00130004000e002b00100000, 128'h10001c000f00000004001e00080007, 128'h1600180007001f000e000000180014, 128'h1d0010000a0018000000000011001a, 128'h1d000a00050026000e00320004000b, 128'h160000000d00090009000e00110025, 128'h500010014003d0012000d0018000d, 128'h8000b00000000000000000004001f, 128'h23000100030000001e000500170019, 128'h130000000e000a0003001700000007, 128'h60011001c0003002f000b00000017, 128'h220004000e00070016000e00000000, 128'h2000000000005001c0013000f0006, 128'h1b0000000b0015000f000b000c000e, 128'h1300150014002400000007000b, 128'h1000150012000b0000000a, 128'h370003002f002f00000014000e000e, 128'h22000b000c00130017000f00000000, 128'h2c00000019000a000000000006001b, 128'h24001e001c00190008003100170023, 128'h16000c00040014000b001300170017, 128'h160000000000000000000c000e0000, 128'h2001b00290005001800250026, 128'h1500370012000b000000000000, 128'h110016000000100000000200130000, 128'h40014000c0015001e00000000001c, 128'h2000270017001300000017, 128'h130017002000310000000000160000, 128'h50000001d0026001d0000000c0004, 128'h2b001400000000000a0010, 128'h120019000b00060028000000000000, 128'h3e000300000000000f00040003, 128'h4600000000000d0000, 128'h300070001000d003d000000000000, 128'h40023002000000000000000000000, 128'h280023000d002600320003000e, 128'h1f000f004d00040021000900030000, 128'h0, 128'h7000500000000002e002600120022, 128'h200000032000a0000000000030000, 128'ha00030000001f0000000600000000, 128'h190000000c0020000d000000000013, 128'h150000000000000032, 128'h17003c0009000d001c0000, 128'h1d0017002e000e0000000000090000, 128'h90000002700000019000500240000, 128'h28000700000000001a000e00180000, 128'h48000a00000015000800000002, 128'h60000002a0000000000080000, 128'h14001f003a000000000000, 128'h7003300170000000c000800000000, 128'h15001f001900040012002400000000, 128'h18000d004e000b0012000200000001, 128'h700000000000000000020, 128'hc001200000000002b000c00040029, 128'h40012000200070000000000040000, 128'h140000000000380000001300000006, 128'h18000e0009000b0000000000000007, 128'h70000000000000005002a, 128'h7001a0003002400180000, 128'h1f0029002000070000001000180000, 128'h9000000140005002c0000, 128'h200000003000000003002800260000, 128'h18000000000023000000000000, 128'h100029000000000000000000000003, 128'hd00140000000d00000000, 128'h3500000000000f000d00000000, 128'h21000c000a00090000001600000000, 128'hd00090035000e0001001500000003, 128'h9000500000002000b000000000024, 128'hf002600000000000000220027, 128'hb000000050005000000040010, 128'h16000a000000340000000c0000000b, 128'h240014000800000000000e00000000, 128'h600000011000000120026, 128'h1001b000a002700040000, 128'h160019000400060000000e00120000, 128'h110022000600190000, 128'h40000004100000000003400140005, 128'h600000000001c00080000001e, 128'h2f001100000003002000000019, 128'h30001002100000000002100000000, 128'hc002800000004001e0000000c001b, 128'h240000000500020000000000030020, 128'h300200005002500000006, 128'he0006000d0001000c00000004001f, 128'hd002200000011002b0002, 128'h40007001b, 128'h18000000000008000f0014000c0005, 128'h80000001200110000001200000000, 128'h1e001a0021001100080000, 128'h1600000003000f000c000d00000000, 128'h190000000900040014000000150000, 128'ha0000000500180008000d00000006, 128'h30000002e0022000f002200000006, 128'h290007000900000025, 128'h240000000a000a0019002600000028, 128'h8000b001e0000000a0015001b0000, 128'h2300130000000a001b0000000a0017, 128'h260000000000240019000000000010, 128'h6000e00130002001e001b000c0015, 128'h20002000000000000000000010009, 128'h1f000b0023001900000022001b0006, 128'h30011000600000000000f, 128'h150000000800000000001200080000, 128'h7000e0015001700000009000c0009, 128'h2000000200020001b00150011002a, 128'h1b0010000000130005000000060000, 128'h80000000e00190018000d000d0002, 128'h220005001600060000000400030026, 128'h1a000000000018002f000100090002, 128'h60000000500040000000500000000, 128'h1f000b0000000a0015000800000016, 128'h13001d000500060003000000140000, 128'h120015000c0008001c000300170010, 128'h700000005001f001c00000001000f, 128'h1a0000001d00080013000e00010016, 128'h700060000000f000d000c000a0018, 128'h200000003001e0005000a00180010, 128'h20019000400020015000100000007, 128'h1200020006000c000600010015000d, 128'h7002100000000001f000600000019, 128'hc0000001100010003001c, 128'h1a000000010000000700060006, 128'h80004000b0011001e001800030010, 128'h1b00030019000c000d000000020000, 128'h5001100210004001a0023000d0007, 128'h1700000006000000080010000f000f, 128'h21000d0012000d000e000900000000, 128'h2600180000001300000014000b0000, 128'h1e00130000002000130002000c0003, 128'h17000b000000190000000a0005000c, 128'hc00000004001200000019000e000e, 128'h9000600000000000e001b000d0023, 128'hc00200003000500390022, 128'h70011001f00100014000000000008, 128'hc0008000d00020008000000010011, 128'h6000b000d000d000e000a00000001, 128'h3000600130000000f0011000c0020, 128'hb00060000000f001c00000008, 128'h1500180020001500000011, 128'h8001a00140001000000140010, 128'hf0028000600150005000c0007, 128'h80000000000030003001f0010000c, 128'h3000e0032000000150000000b, 128'h180032000600050017002000000000, 128'h1300310000000900130002000f0000, 128'h15000a000c0012001600150014, 128'h140009000900120025001c00180003, 128'h300000000000a000b000000000011, 128'h1500190000000c002000200032000e, 128'h60000002c002a000f000000000000, 128'h130000001c0001000b000000000019, 128'h1e0000000800090003001a00000009, 128'h800000005001a0000000000000018, 128'h28000200100019000a000c00070000, 128'h500080000000c000b001700000000, 128'he0000002200080022001600050006, 128'h190009000000000030000000070013, 128'h4001400150005000e0024000e000e, 128'hd00160000001c0003001000050011, 128'h160017000c00100010000a00110000, 128'h200260008000000020000000a0000, 128'hd000a000d0015000f000000000000, 128'h28000c0036001e0041001b0000000c, 128'h20000000000140000000000000029, 128'h15000100000016001000080015000f, 128'hc00190005000b000f000000000000, 128'h18000000000011000a000100030016, 128'h2100040004000f0000001400000011, 128'hd0000001a000000000046, 128'h1500000000002200070016000b0000, 128'h140004002100100000001300070000, 128'h12000000260007000c000700030000, 128'h1d000a001c0000001b000f0010000a, 128'h8000100090000000f00120000000b, 128'h140000000000000007000000000000, 128'h3000a000e001b0000000000000000, 128'h26000000000004000c0000000a, 128'h1800000008000c0005000000000000, 128'h3200010014000f0000000b, 128'h5000a000000070004000100020022, 128'h2000f000000040000001000060012, 128'hd00140005000a0018000100000003, 128'h140000000000160005000000030008, 128'h10000b000000000008000b00000000, 128'h150000000000000000000f, 128'hf0003001300030000, 128'h160004001b00090000000f00140000, 128'h160010000e000900040000, 128'h100090039000000000028000d0000, 128'h3001f0000000e, 128'h21000d000000000006000000000007, 128'h700000005001b0000000000000000, 128'h30012000000000009001000000005, 128'h1f0005000c00110000000000000000, 128'h800130000000b, 128'h60009000400090004000400000011, 128'h80023000500000009000f0000, 128'hc0002000b0001001100020000000c, 128'h140008000000070003000000000006, 128'hb000c000400000005000c00000000, 128'hf0000000d0000000d000a, 128'h30000000000020006001000040003, 128'hb00000008000100170000, 128'h40010001b000700250000, 128'h2003300000000003200000000, 128'ha002600010018, 128'h20002400000000000a001100000000, 128'he000b000900140000002a00000000, 128'hd0000000c00080012000a000c, 128'h130006000000050000000000000013, 128'h180000003500020004, 128'he000600000007000a000600040026, 128'hb00250020000d0009002c000a, 128'h2000000000000000d000400000023, 128'h1a000b00000004000a0000000b000a, 128'h40007000300000003001700000007, 128'h4000000210000000f000d, 128'h500000007001300010001, 128'h3000000000000001a000000100002, 128'hb0021000e00220007, 128'h23002b0000001d00000000, 128'h15000d00250005002f, 128'h40021000000000015002300000022, 128'h2b000c000f00000000002900120000, 128'h2b000e00000022000a0000000d001b, 128'h26000000000013000000000000000d, 128'hd000200000011002f0032001e0010, 128'h50010000000160000000000060020, 128'h130003000c00400003002400350000, 128'h200070006000000000017, 128'h22000000000000000200000005000e, 128'h180000001900190000002600000000, 128'h100000017000e002e001100000021, 128'h160000000a0000000e000700000000, 128'hd00000004000b000e000000070006, 128'h150000001c00140000000f000c000b, 128'ha0013002a003c000000000000, 128'h50000000e001e0000002500000014, 128'h26000100080004001900020000001b, 128'h320015000100080000000000050000, 128'h1a00120019001100100003001d000f, 128'hf0000000000190009000100000007, 128'hb000000160000001c001c000c0011, 128'hd000e0000000c0015000b000d001a, 128'hb0002000c002f00000013002e000b, 128'h20000f000f001a000500000006, 128'h2700000002000c000000000000000e, 128'h12001b000100000015000400000008, 128'he00090018000b00020018, 128'h1600060000000000000000000d, 128'h5000c000e001b001f000d0004000e, 128'h300000015000b00020000000e0009, 128'h30006001f00020031001b00050002, 128'h90000000000000021000d0014, 128'h2800000001001e0020001200060006, 128'h2f00080006001100000006000f0001, 128'h230007001400140000000000030006, 128'h80004001100240007001200020019, 128'hc000c000e0000000a00160016000d, 128'h7000d000000030000000c001c000f, 128'he0010000f001b0009000500330008, 128'h7001c0003000e000a00000006, 128'h9001400120000000e00000000001f, 128'h10000400110007001100160009001a, 128'h2000e000700050010001500150021, 128'hd00180002000a0008000600000000, 128'h150012001f001a000e0013, 128'h2000000280009000a001200120012, 128'h6001900130010001f000b0000000c, 128'h400030000000f000e002500130002, 128'h2900000000001600070000000b0005, 128'h140011000000120010000100150000, 128'h12001c000b00110000000000030002, 128'h10005001d0029000a000900000018, 128'hf00140000001e000d0000000a, 128'h700080000000d00000000001a002d, 128'h170012000700000013001d00230005, 128'h1100210015000100000000000d, 128'h13000000150008000500000000001a, 128'h70006000c0009001c001b00000004, 128'h3000000000000000900130028, 128'h6000000060001001a00020000, 128'h14000000180008000e000e000d000f, 128'h8000000290015002e0008000f0005, 128'hd0020000e001f001d00000000, 128'h10000600000009001e002a00130002, 128'h2c0007000000040012000000000000, 128'h1a000300000023000f000a00170000, 128'h1200110007000b0004000000070008, 128'h80005001a00170001000200000016, 128'h40011001b0000000d00160011000c, 128'h10000c000000100009000400190031, 128'hb00110006001b000c0011000e0003, 128'h6001500080000000900000000000c, 128'h1900010000000a000d000000000024, 128'hc000a000000020018001800000009, 128'h110000000000190005000d0008, 128'ha00000000000d000a000b0000, 128'h120000000600060015000c000d000d, 128'h1800180023000f00090009, 128'h16002e00040008002200040000, 128'h70000000000000000002100110009, 128'h2000000000000d0014000100000000, 128'h9000b00000020000d000000040003, 128'hd000e0006000c00000000000e0008, 128'h12000a0016000f0008000600040014, 128'h8000c000b0000000b000e0017000a, 128'hd00080004000c000a000e0013001a, 128'h13000c000600100016001700020000, 128'ha000a000f00000007000600000010, 128'h19000400000009000b000000000019, 128'hf000d000000080012001800000008, 128'h1000050000000c000c000a000d, 128'hf000000000010000000080000, 128'h80000000a000200160000000a0006, 128'h17001a0015000c0008000a, 128'h1700210005000a002700000002, 128'h40001000000000005002300150008, 128'h2100000003000d000e000200000000, 128'he000a000000220009000000040004, 128'hc000000060009000000010010000b, 128'h16000b0015000d0002000300060013, 128'h8000c00030000000b000700180007, 128'he000d0009000c0005000e0010000d, 128'h1500070004000b0018001000000000, 128'h90000000b0000000300070000000f, 128'h17000800000005000c00000000001c, 128'he000d00000008000d001a0000000b, 128'h1100020000000a000d000a000f, 128'h1000c000000000010000000040000, 128'h90000000e000000160000000b0009, 128'h11001c0011000b000a000a, 128'h1b000b0003000d002700000005, 128'h80002000000030004002400110009, 128'h2f000c0000000d000f000200000002, 128'hd0006000000210000000000000000, 128'hf0002000900080000000000100001, 128'h21001000140016000000000006000d, 128'h5000d000000000010001300180006, 128'h15000a0007000a0005001000120019, 128'h110007001f000c00150006000e0000, 128'hb000000090000000000060000000f, 128'h14000b00000000000d000000000020, 128'h13000c00020007001100190000000b, 128'h11000200000018000d0013000f, 128'h2000e000000000011000900000000, 128'h30000000c000000170000000d000a, 128'hc001b0020000b0029000f, 128'h20017000e0006000d002f00000008, 128'h4000d002a00150019, 128'h2d0012000000030015000000000000, 128'h280002000000140005001300100000, 128'h230007000d000c00060002000c0000, 128'h140010001400130000000500000013, 128'hc000f00000007001e00160009, 128'h1000110000000f0000000500190020, 128'h1500160012001f00130011001a0002, 128'h60007000800000000000000000011, 128'h130005000000100010000000000022, 128'hc000000000000000e001f00000011, 128'hd0000000000160004000f0009, 128'h600000000000b000c00080000, 128'h60000000b0000001e00000013000a, 128'h11000c0017000c00200015, 128'ha00110011001d0019001300000006, 128'h30005002d000c0020, 128'h220009000c00070019000300000000, 128'h2e001300000012000e000b000a000b, 128'h21000f001a002500100000000b0016, 128'hd000e001800190000000f00020016, 128'h8000d0000000b001600110011, 128'h9001e00000018001a000d0020001f, 128'h12000b0005002500040006001f0012, 128'h6001b001200020013000300060006, 128'h23000300000006000c000000000024, 128'h12000e00000000001700170000000f, 128'h13000000000020000800110007, 128'h1b000000000014000300030008, 128'h70000000600110012000300080019, 128'h12001b0008000a000f001a, 128'h1000b001b00060019001e00000004, 128'h2000a00040004002000160008 };

   wire [63:0] airplane4_mp_3_image [1023:0] = { 64'he0011001c0015, 64'h20000900120004, 64'hd00000000, 64'ha0000000f0000, 64'hf001700060000, 64'h13002000160004, 64'h600150028, 64'h230009000a000c, 64'h11001b0018001d, 64'h16000f00380000, 64'h1d0000000c001c, 64'hc000c000c0019, 64'h140008, 64'h3001000030014, 64'h19001200160012, 64'h1c000700130008, 64'h5000a000d0000, 64'h23001b00130005, 64'h12000c0001, 64'h9000800130000, 64'hc001a00080015, 64'h110013, 64'h130009000a0007, 64'h900180020001b, 64'h32000f00000006, 64'h1400000013000e, 64'h1e001700150000, 64'hb00000000, 64'h25000000190000, 64'h13000f00150000, 64'h2000090000000d, 64'h100040006, 64'h1600150003, 64'h8001d00000000, 64'h1b00110013, 64'h230020001b0000, 64'h220010001b001c, 64'h120015000a001a, 64'h1f000a001a0004, 64'h30001c0009000b, 64'h17001300000016, 64'h16000b0000, 64'h17001000000000, 64'h18001300280004, 64'h1000b, 64'hf000000000014, 64'h15000300070000, 64'h16001400080009, 64'he000900030011, 64'hc000100000000, 64'h11001200000011, 64'h9001b0000, 64'h1e00110011, 64'hf0007, 64'h7000e00000000, 64'h160023001a, 64'h14000c00140016, 64'h20000d00000010, 64'h16001500160027, 64'h17000e0015, 64'h60000001c0000, 64'h9000f000c0014, 64'h600290010000e, 64'h5000c00000004, 64'hd0000000d, 64'h110006, 64'h14002700000000, 64'h1b0018, 64'h19001000000000, 64'h8000600000016, 64'h14000b0018, 64'h15001600120009, 64'h2001f001c0015, 64'h70014002f0000, 64'h13000700000034, 64'hf0005002a0025, 64'h13001600070000, 64'hd000100000018, 64'h400280000, 64'h180014001c0000, 64'h9000000150014, 64'he000000110000, 64'ha001400020009, 64'h260000003a0017, 64'h1200000000002c, 64'h6000d000d001f, 64'h150006001e000b, 64'h50000002c0000, 64'h1200000000000d, 64'h1900080000000e, 64'h24001a, 64'h0, 64'h1e000c00210000, 64'h10000d002a0001, 64'hf001000030005, 64'h6000b0000002b, 64'h10, 64'he000f00010017, 64'h1a000000000013, 64'h1f000000090000, 64'hc001e0028, 64'h400030017, 64'h16001c0000000f, 64'h280003000c0002, 64'h100110000000f, 64'h210000000b0000, 64'h11001100120000, 64'h100120000, 64'h500260000000f, 64'h40014, 64'h25002000070000, 64'h18000f00170002, 64'h2a000a0000000c, 64'h2300000000, 64'h2a000000000011, 64'h1000000011, 64'ha001900000012, 64'h1000900000020, 64'h1b000000190000, 64'h150013, 64'h1c001d00000017, 64'h14001100070000, 64'hf000a0000, 64'h1600180000, 64'h1b000a, 64'h900020000, 64'h17000200000017, 64'h6001c00000003, 64'h14000100000017, 64'h700000005001d, 64'h18001a00000001, 64'h13, 64'h15002200000000, 64'h7000800030000, 64'hc0000001f0004, 64'h7000e00210002, 64'hf000800050023, 64'h1500000007000a, 64'h1e0000001f, 64'h1001d0001, 64'h25001200090000, 64'h1a00100000001e, 64'h11001d000b, 64'h1200250000, 64'h700200000, 64'h700000012000d, 64'hb001a00000000, 64'h1a000000300007, 64'h70000001c, 64'h5001300130010, 64'h140000000f0000, 64'h18001800060001, 64'h600000008, 64'h2800000000001a, 64'he00030014002c, 64'hb00160000, 64'h27000500000000, 64'h9000000200000, 64'h1c001600000008, 64'hf00000029, 64'h140000000e, 64'h1500060013, 64'h14000400000009, 64'h70000000d0000, 64'h210004000b, 64'h1c000a0007, 64'h7001100000016, 64'h1100000008000c, 64'h14001400030002, 64'h24000000010017, 64'he0006001b0008, 64'hb000200160000, 64'h4001e000a0000, 64'h100000013, 64'h10001b0004, 64'h5001200000010, 64'h19000d00030003, 64'h1a00000005, 64'h1f00000000001a, 64'h5001500020005, 64'he00150007000f, 64'h2600070000000b, 64'h20000b00060002, 64'h20024, 64'hc001100090002, 64'h13000900000000, 64'hb0000000c0000, 64'h1700070000, 64'h150001, 64'he00110018, 64'h17000f0000000f, 64'h1c001e00000000, 64'h17000800050013, 64'h6001d00000015, 64'h29001000180001, 64'h13000a0008000b, 64'h7002800000010, 64'ha0024000f0000, 64'h2e001f0005, 64'h120000, 64'h9001400000021, 64'hc0006000a0008, 64'h500150027000e, 64'ha0012000e002b, 64'h21000900100010, 64'ha001000090019, 64'h23001c0003, 64'h2100160000, 64'hf00000020001a, 64'h12000000020021, 64'h1900030000, 64'hd00060011000c, 64'h10000000110017, 64'ha0008000c0014, 64'h10001300130010, 64'h1e0000000f000f, 64'hb001300210011, 64'h17000000170011, 64'h24000c0011001b, 64'h1000a00070005, 64'h6000f0011000a, 64'h20000b001d001a, 64'h1c0000001f0013, 64'h3000a002e, 64'h5000500060006, 64'h1c001e00050009, 64'h1500130000000e, 64'ha000100180014, 64'h1000000004, 64'h150009001d0009, 64'h1c002000130013, 64'h50000000d0006, 64'h1a0019000b0000, 64'h19001300000014, 64'h2200140021000e, 64'h230000, 64'he001800000000, 64'ha000000090001, 64'h7000900090012, 64'h9001200180002, 64'h200150010001b, 64'hc001e0002000d, 64'h9000000180022, 64'hb000800230013, 64'h4001400100000, 64'h20000000000016, 64'h1800090001000c, 64'h100026, 64'h19000800060014, 64'hd002100000000, 64'h2100000000000d, 64'h5001100150012, 64'ha000000170013, 64'h8002000090006, 64'h180008000c000e, 64'h18000c000a0000, 64'h3000000080001, 64'h1300010015000c, 64'h900000000, 64'h2000000060000, 64'ha001200160000, 64'h9002200030000, 64'h1e00150010001b, 64'h2f002600140015, 64'h1c001a00000025, 64'h9000000110004, 64'h1000000170008, 64'h6001c0000, 64'h11001a0000, 64'h9000f00060000, 64'h2a000c, 64'h600000000000d, 64'h50000, 64'h12000900190003, 64'h10000800050000, 64'h100000000b0000, 64'h1600000012, 64'h8000000040019, 64'h800000000001d, 64'h14000e000e, 64'h35000500000006, 64'h18000b00130010, 64'h5000000000000, 64'h1200030000, 64'h1a000c00180007, 64'h1c00000008000b, 64'h70024000c0000, 64'hc00060003, 64'hf000e001b, 64'h0, 64'hf0000, 64'h1000f00000000, 64'h30012001f0000, 64'h90017000a0011, 64'ha0000, 64'h8000a00010016, 64'h11000000050007, 64'h700000000, 64'hb001100030000, 64'h1400160013000e, 64'h7000a0004, 64'h15, 64'hc00000000, 64'h2a001a0000001b, 64'h150010000d000a, 64'h0, 64'h2000000000, 64'h12000600010000, 64'he001b000f, 64'h400000000, 64'hd00030000, 64'h2800000020, 64'h70000, 64'hc001700000006, 64'h1400260025000f, 64'h9000a000f0000, 64'hb0000000b0000, 64'h10000000d0000, 64'h2800000000, 64'h14001200030000, 64'h1a0000, 64'h7000700000000, 64'hc0012000f0000, 64'h5000000000000, 64'h18000a00090000, 64'h8000300000009, 64'h2a00020000, 64'h15000100000000, 64'h17002a0000000f, 64'h1d001400030000, 64'h0, 64'h0, 64'ha0000, 64'h1000000000, 64'h200340000, 64'he0000, 64'h22000000000006, 64'hc, 64'h800000000, 64'h12000000000000, 64'h1800000000000d, 64'h6, 64'h2f000000000011, 64'h1b0000000f000c, 64'hf00120000, 64'h6, 64'h9000000150000, 64'h1400000000, 64'h400000000, 64'h3000000030000, 64'hc0004000b0006, 64'h14, 64'h0, 64'h500000000, 64'h200000000, 64'h0, 64'h80000, 64'h2e00000000, 64'h10000000000000, 64'h0, 64'h2000000200000, 64'h0, 64'h15001300000000, 64'h130000, 64'h300000000, 64'h0, 64'h16000400000000, 64'h9000000000000, 64'he000000000007, 64'h0, 64'ha000000190002, 64'h600040000, 64'h200060000, 64'h800000014000a, 64'h16001b0002, 64'h2c0000000d, 64'h10000000000000, 64'h2c001c00060000, 64'h1c001b0001, 64'h50000000a, 64'hc, 64'hd00010000, 64'hd, 64'ha000000000030, 64'h7001c0006, 64'h33000300000000, 64'hb000a002a0000, 64'h1400000000000b, 64'h1e001400230000, 64'h1f00000012, 64'h1500080000, 64'h22000000080000, 64'h800000000001b, 64'h32001400020003, 64'h700000000001c, 64'h0, 64'h0, 64'h800000010, 64'h7000600170000, 64'ha0000000b0000, 64'h3, 64'h0, 64'h600060000000c, 64'hf000000000000, 64'h12000000090003, 64'h60010, 64'h2c00000000000c, 64'h1300330008, 64'h12001f0000, 64'h13, 64'h9000c0000, 64'hf0000001d, 64'hc000000000000, 64'h800130000, 64'h18000000140000, 64'h1e00000000000e, 64'h100004, 64'ha00000000, 64'h60000000a, 64'h0, 64'hd001a, 64'h500000000, 64'he000000000000, 64'hc00000000, 64'h18000000290000, 64'h1b002d00000000, 64'hf00000000, 64'h1e0004, 64'h10017001c, 64'h5001300000003, 64'h2a000100000000, 64'h500000000001e, 64'h900000000, 64'h1001f00000000, 64'h500060000000f, 64'h2400000018, 64'h7000c000c0000, 64'ha0000, 64'h700190000, 64'h200000000, 64'h12000000000001, 64'h3c00000000000e, 64'he000c0025001a, 64'h600000007, 64'h300000019, 64'h0, 64'h1000000000006, 64'h3a, 64'h1c0005001b0000, 64'h1b000c00000000, 64'h2e00210031000f, 64'h14001d00180002, 64'h250000000f0000, 64'hd00100008, 64'ha002000180000, 64'h10000000080000, 64'h3001800080007, 64'h1c000000050000, 64'h19000e001e0022, 64'h0, 64'h1000000010, 64'h28000b000f0007, 64'h20000000f0000, 64'h17001c00220003, 64'h4000400100018, 64'he0000001f0000, 64'h12001700250015, 64'h20000000000000, 64'h600000014000c, 64'h60000000c000e, 64'h160010001b0011, 64'h21000300450013, 64'h90006001c0000, 64'h1f001300250019, 64'h27000000000000, 64'h18, 64'hb000000110000, 64'h210000001d0026, 64'h16000000100016, 64'hd000000030030, 64'h1a000000080003, 64'h6002000000003, 64'h2a0018000f0002, 64'h1e000000000000, 64'h17000000130012, 64'h1100000009, 64'h8002400060000, 64'h1b00000012, 64'h14000700010000, 64'h1500000000, 64'h7000000000002, 64'h120000, 64'h1d002700070018, 64'h70013000f0020, 64'h2500000000001b, 64'hd000800000001, 64'h24, 64'hd001800000007, 64'h2500000017000d, 64'hc0019, 64'h1a002000070000, 64'h11000c00000003, 64'h20015, 64'h500000000000d, 64'h6000a00000000, 64'h2a000200050000, 64'hf0016000f001f, 64'h90016000f, 64'h50000000b0011, 64'h200000006000d, 64'hc000f00150000, 64'h5000b0001002b, 64'h10017000a, 64'h28000000040000, 64'h500000000, 64'hb00000000000f, 64'h6001a00100000, 64'h3003300000000, 64'h9001000010005, 64'h3300220003000a, 64'h1f000f00090010, 64'hb001000090009, 64'hf000700110017, 64'h2200200000, 64'hc, 64'h14000d0000, 64'h200180007, 64'h110007, 64'h0, 64'h140004000f0000, 64'h12000a00150011, 64'h4, 64'h110015000a0007, 64'h1f, 64'h1100000000001c, 64'h6002200240014, 64'h1c00170007000c, 64'hc000000000008, 64'hd000000000000, 64'h110004001c, 64'h23000000050000, 64'h100090000, 64'h2e002a001d0000, 64'h2000120000001f, 64'he00050010, 64'h80003000f, 64'h1b00010003, 64'h1100000000, 64'h10015002b000d, 64'h1f0000000b, 64'h900000010000a, 64'h3001100000000, 64'hc000f00050016, 64'h700000000, 64'h600070001, 64'h1d000400090008, 64'h500050003, 64'hf, 64'h6001700000002, 64'h1000000050014, 64'h17001900000009, 64'h4, 64'h12003100000011, 64'h1002a00000005, 64'h5001f0010, 64'hf0006, 64'hb00120000, 64'h2200000010, 64'h3000b00210000, 64'h1a001800000020, 64'h16001400180000, 64'h2001600120000, 64'h13000000070005, 64'h150000, 64'h16001100000000, 64'h1c00160015, 64'h1a0000001a0002, 64'h1a000000000000, 64'h0, 64'h0, 64'h260000000d0000, 64'h900000000, 64'h1500000000, 64'hf0011000f0000, 64'h8, 64'he000000090000, 64'h70000000a, 64'h500000000, 64'h1a00000000, 64'h17000000040005, 64'h1f0000, 64'hc000500190000, 64'h3000000040000, 64'h12000000000000, 64'h17000d00000010, 64'h7000000000000, 64'h60000, 64'h0, 64'h300000000001c, 64'h17000000120006, 64'h240000, 64'hf0000, 64'h110000001a0000, 64'h0, 64'h2000000040000, 64'h4000000150000, 64'h21000000000001, 64'h15000000000015, 64'h1a, 64'h0, 64'h1f00010000, 64'h0, 64'h200000000f0015, 64'h2b00000000, 64'h2000000000, 64'h0, 64'ha000000030000, 64'hb00000000, 64'h0, 64'hf0000, 64'h230000, 64'h11, 64'h17000000000008, 64'h12000000000000, 64'h0, 64'h0, 64'hc00120000000a, 64'h0, 64'h8000d0000, 64'hd0000000a0000, 64'h0, 64'h1100000010, 64'hf00000000, 64'h18000900000007, 64'h12001c0023000b, 64'h9000f000b0010, 64'h1b, 64'h0, 64'h1c000b00000018, 64'h400000037, 64'h28000d001e0014, 64'h2000000000000, 64'h400000000, 64'h700000000, 64'h33000000060000, 64'h0, 64'h0, 64'h15000f00110000, 64'h13000a00000025, 64'h18000000160000, 64'h400000013, 64'h0, 64'hb001300000000, 64'h23000000000001, 64'hd000000100002, 64'h140002000a0000, 64'h0, 64'hd000c00110000, 64'h4000500180007, 64'h0, 64'h700130000000e, 64'h0, 64'h11000000000016, 64'h3d0007, 64'h18000000160000, 64'h180000, 64'hc0000000e0000, 64'h1800000017, 64'h12000000040000, 64'h2c0000, 64'h17000000000000, 64'h7000000000004, 64'h24000b, 64'h0, 64'h4000c00040000, 64'ha000800000000, 64'hb00000031001b, 64'h1b00000000, 64'h600000000, 64'h200000000, 64'h150000, 64'h700000000, 64'h0, 64'h0, 64'h400080019, 64'h7, 64'h42000000000000, 64'h5000000000018, 64'he, 64'h0, 64'h2, 64'h0, 64'h700030000, 64'h50000, 64'h1700000006, 64'h0, 64'h16000000000000, 64'h11000000000000, 64'h1e001400000016, 64'h2000a0000, 64'h0, 64'h0, 64'hd00000000000d, 64'h5000000000036, 64'h24000200000000, 64'hf000a000d, 64'h1300300012001c, 64'h18001600110016, 64'h1400000010000e, 64'h1200000008, 64'he000100060008, 64'hc001b000b0013, 64'h1c000b0000000d, 64'h15000a, 64'hc00000000001a, 64'h12000000000000, 64'h2001100120012, 64'h2b000000130000, 64'hc0000, 64'h6000d00000013, 64'h12000d000b000b, 64'h13000000190019, 64'h170001000e0028, 64'hc, 64'h100090005000c, 64'h50007000c0007, 64'h9000e0000000d, 64'hf000200350002, 64'hb000000000002, 64'h7001500160015, 64'h16000000050000, 64'h400020000000f, 64'ha00140023000b, 64'h1c0006001d0018, 64'h11001600070007, 64'h12, 64'h1100000012, 64'h40000000d, 64'h16000c00150019, 64'h2900000000000a, 64'h11000000130024, 64'h1800000016, 64'h600090000, 64'ha00060002001b, 64'h1200120003, 64'h2, 64'h6001100070000, 64'h2000000110000, 64'h13000e0000000a, 64'h1700090013, 64'h1f000000000000, 64'h29000c0000000b, 64'h500060002001c, 64'h18001300000000, 64'h1b00100014000a, 64'hd0000, 64'h12000e00160001, 64'h9000500000016, 64'h1600130010, 64'h3, 64'hf001b00000000, 64'h10000000140000, 64'h20015000d0008, 64'h5001c0005, 64'h600000002000f, 64'hd000d00120000, 64'h13000000000006, 64'h1a0000000c0010, 64'he000d00210024, 64'h1c001900120014, 64'h1f000d0000001d, 64'h6001e00020010, 64'h8000e00180019, 64'h190009000e, 64'h1300050000001a, 64'h2200250005001a, 64'h150004000e0008, 64'h1c000000080000, 64'h200050012000a, 64'h7001000040000, 64'h1b000d0010, 64'h6000e000e000c, 64'h12000b00140017, 64'h600000000001c, 64'ha0000001c, 64'h24000c000e0000, 64'h16000d00020012, 64'h1000300000011, 64'hf001500210000, 64'h190000000d0000, 64'h8001400010015, 64'h6001900170004, 64'h50015001a, 64'h15001400040005, 64'h9001400000008, 64'h120019001d, 64'h1200230012000a, 64'h1a001100000007, 64'h190011001f000a, 64'he00140003000a, 64'hf001b0015001a, 64'h170000000d0003, 64'h3001b00140000, 64'h1e00000001, 64'h15000b001b0013, 64'h20008, 64'hb0010000a000a, 64'h900180007, 64'h2001600180025, 64'h8001200000009, 64'h1200040005, 64'h19000900140012, 64'h1700140008, 64'he0016000f0009, 64'h10000000000002, 64'hd000800000012, 64'hb000f000d0003, 64'h80000000d000e, 64'h90029000f000a, 64'h10001b00040009, 64'h40002001d0010, 64'h12000f00190000, 64'h6000c00070006, 64'h8001a000a000d, 64'h9001500190005, 64'h18001400070010, 64'hd001d002a0009, 64'h150024001a0000, 64'hf00090007000e, 64'hf00170000, 64'h1c002000050002, 64'h8000800110015, 64'h1a0012000e0022, 64'h12002300000008, 64'h1c000700050022, 64'h2a00030000, 64'ha0000001d0010, 64'h9000a0000, 64'h16000000000000, 64'h190017001b000c, 64'h10000500000000, 64'h130000000a0005, 64'h7000000080007, 64'hc000100040006, 64'h5000a00000014, 64'h26000000040000, 64'h10000000010015, 64'h17000000020017, 64'h60000000f, 64'h2b001000000000, 64'h1b00000011000a, 64'h60000, 64'h1200180000, 64'ha000000150000, 64'h17000a0001, 64'h3001c0000, 64'h4000000200003, 64'h10001c00080011, 64'h3000000000000, 64'h6001d000f000b, 64'h7000f0000000e, 64'hc0000000c0000, 64'h180010001a0000, 64'h6000600000000, 64'h21001000050015, 64'hf000000000000, 64'h1d001900170007, 64'h600000006, 64'h13000c00100001, 64'h600000000, 64'h1800040001, 64'hc000d, 64'h80004000f0008, 64'h1000000000008, 64'h10000d0000000b, 64'h120010, 64'h1800050000, 64'h2000400080012, 64'h140000000c0000, 64'h1200000000000e, 64'h9000a00000006, 64'h110000, 64'h2000400080003, 64'h19000d00040001, 64'h10000800020014, 64'hd0000, 64'h3000000000003, 64'h800000000, 64'h4001900060000, 64'h300090006000c, 64'h60018000c0000, 64'h1a00180000, 64'h17000400000006, 64'h110000, 64'h18001000000000, 64'h80007000a000f, 64'h1a001c00250000, 64'h900000010, 64'h1c00180009000a, 64'h1b00020000, 64'h230004, 64'hf00080006, 64'h18001200070004, 64'hf001400130002, 64'h1200110000000a, 64'h110004, 64'hf0004000f0000, 64'h80004, 64'h400150008000f, 64'h310000000b0013, 64'h2000000000020, 64'h11000000000007, 64'h80000000a, 64'h15000900010000, 64'h12000000140000, 64'h0, 64'hb0008001a0000, 64'h10000000000000, 64'h1000080014, 64'h40009000f0000, 64'h2000000100002, 64'h5002500070000, 64'h1000900000000, 64'hd003500000000, 64'h18001900060018, 64'h1800000008000c, 64'h900150008000a, 64'h600000007000e, 64'h1d00070000000f, 64'h7000000060000, 64'h1400090011000b, 64'h1100000005, 64'h9001700180000, 64'h10018000b0004, 64'h0, 64'h20000000b0015, 64'h13000000150005, 64'h0, 64'h8001100000000, 64'h20013, 64'he00140000, 64'h100006000f, 64'hc0000000b0000, 64'h11000f00000010, 64'he000600000017, 64'h1, 64'h1400060000, 64'h13000600170000, 64'he00080006000d, 64'h5000000150000, 64'h1e00070000, 64'h500000000, 64'h1900070000, 64'h50000000e001f, 64'h1b00170000, 64'h1000140000, 64'h9000a0011000d, 64'h5000300040000, 64'h900000004, 64'h1e00000007000d, 64'hf00100013001b, 64'h1d00010004, 64'h13001a00080018, 64'h18001700010014, 64'h2000000140020, 64'h14000800100009, 64'h12001500080000, 64'h1500100010001d, 64'h1c000900000000, 64'h600000011001b, 64'hb000c00170011, 64'h900080003000b, 64'h140012001a, 64'h1a000f000b0018, 64'ha000500140023, 64'h100019000a0017, 64'h7001400040019, 64'h19001500020008, 64'h50007000b0006, 64'h500080016, 64'h1d000100160013, 64'h10000d001a0000, 64'h1a00040006, 64'h160007000e0005, 64'ha000d00190000, 64'h1000140008000a, 64'h8000c00130000, 64'h12000000040003, 64'h6002400190011, 64'h170002000a000f, 64'hf000c00190003, 64'h16000700110012, 64'h1100000011000c, 64'ha0003000e0000, 64'h12000c0009000e, 64'h7001200000017, 64'h600000014000a, 64'h20015000a, 64'h110015000d0011, 64'hd000000140000, 64'h40015000e, 64'hf00000002000e, 64'h600110010000e, 64'h7000000150005, 64'hc001f00180000, 64'h14002500180001, 64'hb000000020000, 64'hb00000015000a, 64'h1f00000001000e, 64'hc001d0010001c, 64'h1400170024000c, 64'hf001a00180002, 64'h10000000190018, 64'h15000900150004, 64'h40019000c0008, 64'h9000b00020000, 64'he001a000d0000, 64'h7000d0013001d, 64'h7001e00170000, 64'h5000e001a000c, 64'h12, 64'h14001b0000, 64'h10000f00000010, 64'hd001200100000 };

   wire [15:0] airplane4_fc_1024_preBN_image [1023:0] = { 16'hf9a1, 16'hfe09, 16'hfb75, 16'hffca, 16'h5d, 16'hd9, 16'h117, 16'hfda8, 16'hfcd2, 16'hfb90, 16'h101, 16'h281, 16'hfebe, 16'ha5, 16'hfca7, 16'hfcec, 16'hfc02, 16'hfcd8, 16'hfd86, 16'hfd71, 16'h110, 16'h4dc, 16'hfe5d, 16'hb3, 16'hfe03, 16'hfeda, 16'hfb4d, 16'h307, 16'h201, 16'hfbc4, 16'hff3c, 16'hca, 16'h180, 16'hfeaa, 16'h340, 16'hc4, 16'hfd9f, 16'h11e, 16'hffbb, 16'h4d8, 16'hfebc, 16'h29, 16'hfe01, 16'he4, 16'hff3c, 16'hfea6, 16'hfcf0, 16'hfed0, 16'h13f, 16'h3a, 16'h5ea, 16'hfdbc, 16'h14d, 16'hff51, 16'hfe85, 16'hfe5b, 16'hf918, 16'hfe34, 16'h101, 16'h3d5, 16'h121, 16'hfc8f, 16'hfd9b, 16'hffab, 16'hfe41, 16'h51, 16'hfa56, 16'h53, 16'hff25, 16'hfcbf, 16'h43, 16'h13, 16'h191, 16'hfe73, 16'hfe88, 16'h1d0, 16'hffdc, 16'h1fb, 16'h17f, 16'h1df, 16'hfce2, 16'h24b, 16'h1fd, 16'hff64, 16'hffd3, 16'h3f, 16'hfdf4, 16'hfee1, 16'hfe75, 16'h238, 16'h86, 16'h4a2, 16'hfdc3, 16'h323, 16'hfc71, 16'hfb87, 16'hfe30, 16'hfc3a, 16'h31b, 16'hff5a, 16'hfd85, 16'hff3d, 16'hffa0, 16'hfcc1, 16'h64b, 16'h16c, 16'h226, 16'hfcf4, 16'hfda5, 16'h13d, 16'h266, 16'h2, 16'h1a, 16'hfaae, 16'hffe2, 16'h17f, 16'hfdfb, 16'hfaed, 16'hffd3, 16'hb2, 16'hfed7, 16'hfd8b, 16'hfebf, 16'h41b, 16'h32, 16'h99, 16'hffdd, 16'h308, 16'hfd50, 16'hff7e, 16'hffc8, 16'hfbfb, 16'hff12, 16'h24e, 16'hbb, 16'hfcd9, 16'hffbb, 16'hfe4d, 16'hfe5a, 16'hfda9, 16'hfe50, 16'he2, 16'hff5f, 16'hfe8d, 16'hfea2, 16'hffcd, 16'hfe9b, 16'hff93, 16'hfead, 16'h168, 16'hfec6, 16'hfe1b, 16'hfbc7, 16'hffef, 16'h65, 16'hf907, 16'h4f4, 16'h26d, 16'hfebb, 16'hff3b, 16'hfeba, 16'hfbcb, 16'h154, 16'hfdeb, 16'h5d, 16'h140, 16'h1f5, 16'h1ea, 16'hfff4, 16'hfd33, 16'hfe99, 16'hfb79, 16'h203, 16'hfda4, 16'hff1a, 16'hfe95, 16'hff3b, 16'hfe08, 16'hff07, 16'hfbd7, 16'h1ee, 16'hfcc4, 16'hff4f, 16'hfd63, 16'hfda2, 16'hfc9a, 16'hff2f, 16'hfd60, 16'h71, 16'hfdbc, 16'hfd50, 16'hfe6b, 16'hfd17, 16'hfe8a, 16'hffde, 16'h131, 16'hff86, 16'hfe9e, 16'hfdcf, 16'hfedb, 16'h245, 16'hffb1, 16'hfc0b, 16'hfcd7, 16'hfe8b, 16'h6f, 16'hfe40, 16'hff49, 16'hfe74, 16'hffb7, 16'h112, 16'hfdba, 16'h323, 16'hff4e, 16'hff50, 16'hfcb3, 16'hfe56, 16'hff73, 16'h23, 16'hff92, 16'hfff3, 16'hfe09, 16'hff4b, 16'hfd89, 16'hfffd, 16'hff53, 16'h281, 16'h135, 16'hfee7, 16'hfacf, 16'hff51, 16'h15d, 16'hfceb, 16'h2bb, 16'hfa96, 16'hfeba, 16'h15e, 16'hc2, 16'h42f, 16'h50a, 16'h345, 16'hfbae, 16'hff05, 16'hfdc7, 16'hfc5f, 16'hfe85, 16'hfd8f, 16'hfffc, 16'hfd5c, 16'h1a0, 16'hfe25, 16'h461, 16'h36, 16'h166, 16'hfe0f, 16'hff66, 16'hfd4b, 16'hffb7, 16'hbc, 16'hfe28, 16'hff76, 16'hfe04, 16'hfd20, 16'hff3f, 16'h299, 16'hfea3, 16'hfdc2, 16'hfaf2, 16'hfcec, 16'hfebd, 16'hfafb, 16'hf8, 16'h3a3, 16'hff75, 16'hfdcc, 16'hfeb0, 16'hfee4, 16'h209, 16'hfd95, 16'h3e7, 16'hff99, 16'hfdbf, 16'h61, 16'h282, 16'hfff1, 16'h2a9, 16'hfe51, 16'hfd13, 16'hfd7a, 16'hfb73, 16'hfb18, 16'hffef, 16'h2b5, 16'hfd07, 16'hff71, 16'hffcb, 16'hfd33, 16'h145, 16'hfcce, 16'h6c0, 16'hfbb7, 16'hffce, 16'hfec3, 16'hfdee, 16'hfd5b, 16'h259, 16'hfc9a, 16'hfc32, 16'hfdab, 16'hfbe8, 16'hfb3b, 16'hfe10, 16'h3e3, 16'hfd40, 16'hfe56, 16'hfeee, 16'hff36, 16'h112, 16'h2c1, 16'hfd2d, 16'hff43, 16'hfe8e, 16'hff3f, 16'hf9cd, 16'hfeda, 16'hfdd0, 16'h9f, 16'hfbc6, 16'h172, 16'hca, 16'hfe74, 16'h1bb, 16'hfba2, 16'hfc28, 16'hfc34, 16'h465, 16'h138, 16'hff0f, 16'h11b, 16'hfdcd, 16'h39e, 16'hfcef, 16'hfd84, 16'hfef4, 16'hfd2a, 16'hffc4, 16'h565, 16'hff67, 16'hfdc1, 16'h3a3, 16'h137, 16'h53, 16'hfc52, 16'hfe6f, 16'h126, 16'hff73, 16'hfd22, 16'hfc21, 16'h5ce, 16'h43, 16'hfd2e, 16'h63, 16'hce, 16'hfa05, 16'h104, 16'h25e, 16'h5e, 16'hfb56, 16'h1e, 16'h76, 16'hfdbf, 16'h280, 16'h1ab, 16'hff7b, 16'hff00, 16'hfcdf, 16'hfee6, 16'hff9c, 16'hfd04, 16'hfee5, 16'hff47, 16'h349, 16'hfd67, 16'h21f, 16'hfb82, 16'hfe87, 16'hff7f, 16'h2ec, 16'hfe92, 16'hfb52, 16'h20, 16'h50a, 16'h134, 16'hfec9, 16'hfe75, 16'hfe17, 16'h230, 16'h118, 16'hfefc, 16'h175, 16'h10d, 16'hfff0, 16'hff16, 16'h385, 16'hfbf9, 16'hfcc0, 16'hfddc, 16'hfec4, 16'h189, 16'hfd32, 16'hfc6f, 16'h2d4, 16'hfec0, 16'h176, 16'hfdae, 16'hffbe, 16'h3a6, 16'h12, 16'h21d, 16'hfe75, 16'hfc2f, 16'h2f8, 16'h10d, 16'h215, 16'hf, 16'hfd1b, 16'h1df, 16'hfa, 16'hfae2, 16'hfc81, 16'hfdc7, 16'hfda1, 16'hffb2, 16'hfbf7, 16'h38, 16'h327, 16'hfdd1, 16'h1f, 16'h128, 16'hfbbe, 16'h1d5, 16'hffa7, 16'hffcc, 16'hffee, 16'hfb3d, 16'hfd0f, 16'hffc9, 16'h138, 16'hfed5, 16'h3c3, 16'h288, 16'h108, 16'hfdc3, 16'hfb1f, 16'hff7d, 16'hfc0f, 16'hfe6c, 16'hfc13, 16'hffdf, 16'h5cb, 16'h1ef, 16'hfd48, 16'h2a5, 16'hfcef, 16'hffca, 16'hfbaf, 16'hf8b9, 16'hfeb0, 16'hff92, 16'hfe66, 16'h419, 16'hfeaa, 16'hff8b, 16'hffd5, 16'hff31, 16'h25, 16'hfe30, 16'h21, 16'hfea7, 16'h513, 16'h3d8, 16'hff09, 16'h244, 16'hfe2f, 16'hc7, 16'hfb7b, 16'h58, 16'h402, 16'hfe96, 16'hfa93, 16'h2e, 16'hfa81, 16'hfdde, 16'hfecd, 16'h4e6, 16'hfe73, 16'hff21, 16'hfce4, 16'hfdb8, 16'h584, 16'hffb4, 16'h8d, 16'h306, 16'hfc85, 16'hfe81, 16'hfff6, 16'hfca0, 16'hfd92, 16'hff18, 16'h48b, 16'hfbb2, 16'hfdb7, 16'hfe68, 16'hfe99, 16'hfe72, 16'hfce7, 16'hfde4, 16'he2, 16'h6f, 16'hfec3, 16'ha5, 16'hfe98, 16'hfa29, 16'h40c, 16'hfdd1, 16'he, 16'hfdc4, 16'hfdcf, 16'h59d, 16'hfece, 16'hfde5, 16'h79, 16'h12c, 16'hff03, 16'hfc5a, 16'hfef6, 16'hfa7e, 16'h26e, 16'h21d, 16'hff44, 16'hfbc8, 16'hfead, 16'hfda3, 16'h121, 16'hfd70, 16'h37, 16'hfc3f, 16'h32, 16'hfe94, 16'h176, 16'h8f, 16'hfd74, 16'hf8ec, 16'hfcff, 16'hffcc, 16'h26, 16'h2ca, 16'h18b, 16'h85, 16'h29e, 16'hffb6, 16'hfd0f, 16'hfc6c, 16'hfe99, 16'hfe28, 16'hfe37, 16'hfc54, 16'hfd79, 16'h461, 16'h2a9, 16'hfd5b, 16'hfd68, 16'hff14, 16'h714, 16'hfe20, 16'h9f, 16'hfd8b, 16'hb7, 16'hffe4, 16'hfe6d, 16'h7f, 16'hffe1, 16'hf98f, 16'hfe6c, 16'h2c9, 16'hffa4, 16'hfc47, 16'h543, 16'h191, 16'h469, 16'hfd75, 16'h273, 16'hfe5d, 16'hfc4d, 16'h107, 16'hfdbc, 16'hfd84, 16'hfd2f, 16'hfcab, 16'h2e3, 16'h1f0, 16'hfd7a, 16'hfcad, 16'h1d3, 16'hffd8, 16'hfe8f, 16'hfe8a, 16'h2e3, 16'hfccb, 16'hc2, 16'hfe7e, 16'hfb38, 16'hff1e, 16'hfff4, 16'hff84, 16'hfe66, 16'hfd6a, 16'hf6, 16'haf, 16'hff78, 16'hfc17, 16'hfc2d, 16'h36, 16'hfcde, 16'hfd4b, 16'hffd0, 16'h262, 16'h11e, 16'h23, 16'he7, 16'hff7a, 16'h1f4, 16'hfec9, 16'h155, 16'hfc8f, 16'hfda2, 16'h25, 16'h157, 16'hff66, 16'hfcba, 16'hfda1, 16'hfc7f, 16'hfedd, 16'h1fe, 16'hff60, 16'h219, 16'h6d1, 16'hff52, 16'h2f8, 16'hfe6e, 16'hfdab, 16'hfcc1, 16'hf934, 16'hff26, 16'hfee6, 16'hff64, 16'hfdae, 16'hfdc2, 16'h24b, 16'hfd26, 16'h3e5, 16'hfe9e, 16'hff8f, 16'h14f, 16'hfc70, 16'h2f1, 16'h15e, 16'h33e, 16'h153, 16'hfdd4, 16'hfb69, 16'h218, 16'hfc56, 16'hfd92, 16'hfd4c, 16'hff7e, 16'h280, 16'hfcc6, 16'h1d9, 16'hfd35, 16'hfe86, 16'hfdde, 16'hfc8d, 16'hf944, 16'hfb31, 16'h95, 16'hfe8b, 16'h13b, 16'hfefc, 16'h211, 16'hfc66, 16'hf963, 16'h3a4, 16'hc5, 16'hfb16, 16'hff22, 16'h4a3, 16'h14c, 16'hfe72, 16'hfd01, 16'hfdb1, 16'h2fc, 16'ha2, 16'hffb8, 16'hfdd3, 16'h2b0, 16'h158, 16'hfbf7, 16'h19f, 16'h8f, 16'hfef8, 16'hc5, 16'hffc0, 16'h30, 16'hfe11, 16'h10c, 16'h27f, 16'hff41, 16'hfb7f, 16'h11d, 16'hfe17, 16'h2f9, 16'hfde0, 16'h294, 16'hfc44, 16'hfec7, 16'hfefa, 16'hff08, 16'h112, 16'h1e, 16'hfdbe, 16'h1e1, 16'h3e, 16'hff0f, 16'hffa5, 16'hfc39, 16'hfba4, 16'hfe3d, 16'h37d, 16'hfc79, 16'hff99, 16'hfd9b, 16'hfd02, 16'hfea2, 16'hfe24, 16'hfd4b, 16'h1b, 16'hfd27, 16'h7f, 16'hffd1, 16'h2e, 16'hff81, 16'h401, 16'h2b0, 16'hfd78, 16'hff11, 16'hff7a, 16'hfdd6, 16'hfd70, 16'h84, 16'hfe20, 16'hfb7f, 16'hfd02, 16'hfda0, 16'hfdae, 16'h110, 16'h18b, 16'hfd27, 16'hfcd6, 16'h4, 16'hfce0, 16'hff8e, 16'h73, 16'hfc47, 16'hfd77, 16'hff59, 16'h2b3, 16'hfee8, 16'h1bc, 16'hc2, 16'h23d, 16'h248, 16'h1ae, 16'h260, 16'hf7e9, 16'h3bf, 16'hfbf1, 16'hfef8, 16'hff57, 16'h1ed, 16'h162, 16'h1b1, 16'h5e, 16'hfe5b, 16'hffc3, 16'h43, 16'hff42, 16'hfdbf, 16'h1b8, 16'hfdb8, 16'h2bf, 16'hf7, 16'h19, 16'hfe47, 16'h108, 16'hfd7e, 16'hfe4e, 16'hfec1, 16'hffe3, 16'h2fb, 16'hfeff, 16'h7a, 16'hff63, 16'hfed9, 16'h90, 16'hfbde, 16'hfc60, 16'h33f, 16'hfee4, 16'hff4c, 16'h1f7, 16'hfe81, 16'hfd0f, 16'h1a7, 16'h86, 16'hff64, 16'h4eb, 16'hfec4, 16'h7c, 16'h315, 16'hd3, 16'h42a, 16'hfcbe, 16'hffa4, 16'hfe35, 16'hfdc9, 16'hffdc, 16'hff71, 16'h15b, 16'h2aa, 16'h17, 16'hfe33, 16'h18f, 16'h29b, 16'hfd03, 16'hfb09, 16'hfeed, 16'h353, 16'h6f, 16'h2f, 16'ha1, 16'h1a9, 16'hfec1, 16'h314, 16'hfd19, 16'hcd, 16'hfd84, 16'hfdcb, 16'hff3e, 16'h1c8, 16'hfd5d, 16'hf9, 16'hffe9, 16'h28b, 16'h362, 16'hfeed, 16'hbe, 16'hffd6, 16'h1e, 16'h3ba, 16'h159, 16'hfdb9, 16'hb5, 16'hfe8f, 16'hff5d, 16'h99, 16'hffd2, 16'h20d, 16'hfe04, 16'hff81, 16'hfee5, 16'hfc6e, 16'hc0, 16'hf9dd, 16'h1, 16'hfbf7, 16'hfe05, 16'hfacb, 16'hfbaa, 16'h2d0, 16'hfcf7, 16'hff20, 16'hff3b, 16'h15b, 16'hfedb, 16'hfdd8, 16'hfdce, 16'h96, 16'hd2, 16'hfea8, 16'h23b, 16'h21f, 16'hff3e, 16'hff8d, 16'h1f2, 16'hfa50, 16'hff0d, 16'h201, 16'h18, 16'hfe96, 16'hfbf9, 16'hfdff, 16'hfd6e, 16'hff61, 16'h32b, 16'hff1a, 16'h169, 16'hff42, 16'hfb4e, 16'hff91, 16'hfdeb, 16'hfd1d, 16'hff23, 16'h705, 16'hf904, 16'hffdc, 16'hfe56, 16'hd0, 16'hfee5, 16'hc4, 16'hfe9b, 16'hfc, 16'hffed, 16'hfdce, 16'hfe83, 16'hfe20, 16'hdd, 16'hfc17, 16'h155, 16'h2da, 16'hf9f7, 16'hfb12, 16'hfd6b, 16'h423, 16'hfc03, 16'hffa7, 16'h3f, 16'hfe45, 16'h2c1, 16'h34c, 16'hff1d, 16'hfec7, 16'hfe11, 16'hfbf0, 16'hfda5, 16'h376, 16'hfe54, 16'h4f, 16'h617, 16'hfa36, 16'hfd9d, 16'hfc18, 16'hf4, 16'h327, 16'hff12, 16'h17, 16'hfd9b, 16'hfd35, 16'h3e0, 16'hfb68, 16'hff71, 16'hffbb, 16'hff62, 16'hb3, 16'hff29, 16'hfdc8, 16'hfad4, 16'hfe93, 16'hfef0, 16'hfead, 16'h161, 16'hfdc0, 16'hff9d, 16'hff4a, 16'hfe0e, 16'hfc1b, 16'hfb54, 16'hf8ea, 16'hff21, 16'h127, 16'hfc00, 16'h88, 16'hfaf0, 16'hae, 16'h15d, 16'hfebd, 16'h285, 16'h290, 16'hff37, 16'hff69, 16'hff4b, 16'hfda3, 16'h1fd, 16'hfea5, 16'hfbab, 16'h1b2, 16'hfc20, 16'hfac5, 16'hff48, 16'h74, 16'hfcdc, 16'hfc21, 16'hfe21, 16'hfe88, 16'hfff0, 16'hfedc, 16'h32, 16'hfe05, 16'hffbd, 16'hffc3, 16'hfa23, 16'h2fc, 16'hfcff, 16'ha5 };
   
   reg         clock;
   reg 	       reset;
   wire        rdy_in;
   reg 	       vld_in;
   wire [15:0] bits_in_0;
   wire [15:0] bits_in_1;
   wire [15:0] bits_in_2;
   reg 	       rdy_out;
   wire        vld_out;
   wire [15:0] bits_out_0;
   /*
   wire [15:0] bits_out_1;
   wire [15:0] bits_out_2;
   wire [15:0] bits_out_3;
   wire [15:0] bits_out_4;
   wire [15:0] bits_out_5;
   wire [15:0] bits_out_6;
   wire [15:0] bits_out_7;
    */

   reg 	       start_data;
   reg [9:0]   img_cntr;
   reg [9:0]   out_cntr;
   wire        bits_out_0_correct; /*,
	       bits_out_1_correct,
	       bits_out_2_correct,
	       bits_out_3_correct,
	       bits_out_4_correct,
	       bits_out_5_correct,
	       bits_out_6_correct,
	       bits_out_7_correct; */
   wire [47:0] curr_pixel;
   assign curr_pixel = airplane4_image[img_cntr];

   assign bits_in_0 = curr_pixel[15:0];
   assign bits_in_1 = curr_pixel[31:16];
   assign bits_in_2 = curr_pixel[47:32];
   assign bits_out_0_correct = ( bits_out_0 == airplane4_fc_1024_preBN_image[out_cntr][15:0] );
   /*
   assign bits_out_0_correct = ( bits_out_0 == airplane4_mp_3_image[out_cntr][15:0] );
   assign bits_out_1_correct = ( bits_out_1 == airplane4_mp_3_image[out_cntr][31:16] );
   assign bits_out_2_correct = ( bits_out_2 == airplane4_mp_3_image[out_cntr][47:32] );
   assign bits_out_3_correct = ( bits_out_3 == airplane4_mp_3_image[out_cntr][63:48] );
   assign bits_out_4_correct = ( bits_out_4 == airplane4_mp_2_image[out_cntr][79:64] );
   assign bits_out_5_correct = ( bits_out_5 == airplane4_mp_2_image[out_cntr][95:80] );
   assign bits_out_6_correct = ( bits_out_6 == airplane4_mp_2_image[out_cntr][111:96] );
   assign bits_out_7_correct = ( bits_out_7 == airplane4_mp_2_image[out_cntr][127:112] );
    */
   
   /* Instantiation of top level design */
   AWSVggWrapper
     dut (
	  .clock( clock ),
	  .reset( reset ),
	  .io_dataIn_ready( rdy_in ),
	  .io_dataIn_valid( vld_in ),
	  .io_dataIn_bits_0( bits_in_0 ),
	  .io_dataIn_bits_1( bits_in_1 ),
	  .io_dataIn_bits_2( bits_in_2 ),
	  .io_dataOut_ready( rdy_out ),
	  .io_dataOut_valid( vld_out ),
	  .io_dataOut_bits_0( bits_out_0 )
	  /*
	  .io_dataOut_bits_1( bits_out_1 ),
	  .io_dataOut_bits_2( bits_out_2 ),
	  .io_dataOut_bits_3( bits_out_3 ),
	  .io_dataOut_bits_4( bits_out_4 ),
	  .io_dataOut_bits_5( bits_out_5 ),
	  .io_dataOut_bits_6( bits_out_6 ),
	  .io_dataOut_bits_7( bits_out_7 )
	   */
	  );

/* Add stimulus here */
always #2 clock = ~clock;

always @(posedge clock)
  begin
     if ( start_data & vld_in & rdy_in )
       begin
	  img_cntr <= img_cntr + 1'h1;
       end
     if ( vld_out )
       begin
	  out_cntr <= out_cntr + 1'h1;
	  if ( !bits_out_0_correct )
	    begin
	       $display("Bits 0 out is incorrect");   
	    end
	  /*
	  if ( !bits_out_1_correct )
	    begin
	       $display("Bits 1 out is incorrect");   
	    end
	  if ( !bits_out_2_correct )
	    begin
	       $display("Bits 2 out is incorrect");   
	    end
	  if ( !bits_out_3_correct )
	    begin
	       $display("Bits 3 out is incorrect");   
	    end
	  if ( !bits_out_4_correct )
	    begin
	       $display("Bits 4 out is incorrect");   
	    end
	  if ( !bits_out_5_correct )
	    begin
	       $display("Bits 5 out is incorrect");   
	    end
	  if ( !bits_out_6_correct )
	    begin
	       $display("Bits 6 out is incorrect");   
	    end
	  if ( !bits_out_7_correct )
	    begin
	       $display("Bits 7 out is incorrect");   
	    end
	   */
       end
  end
initial begin
$timeformat(-9,3,"ns",12);
end
initial begin
   clock = 0;
   reset = 1;
   vld_in = 0;
   rdy_out = 1;
   start_data = 0;
   img_cntr = 0;
   out_cntr = 0;
   #32
   reset = 0;
   #32
   // start sending data
   start_data = 1;
   while ( 1 == 1 )
     begin
	vld_in = 1; // $urandom % 2;
	#4;
     end
end

endmodule // aws_vgg_testbench
